magic
tech sky130A
magscale 1 2
timestamp 1762640459
<< metal1 >>
rect -100 100 100 157
rect -100 -157 100 -100
<< rmetal1 >>
rect -100 -100 100 100
<< labels >>
rlabel metal1 0 140 0 140 0 R1
port 1 nsew
rlabel metal1 0 -140 0 -140 0 R2
port 2 nsew
<< properties >>
string gencell sky130_fd_pr__res_generic_m1
string library sky130
string parameters w 1 l 1 m 1 nx 1 wmin 0.14 lmin 0.14 class resistor rho 0.125 val 125.0m dummy 0 dw 0.0 term 0.0 roverlap 0 doports 1
<< end >>
