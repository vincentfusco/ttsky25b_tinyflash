** sch_path: /home/bmott/ttsky25b_tinyflash/xsch/ip/top/tt_um_flash_adc/tt_um_3bit_flash_adc.sch
.subckt tt_um_3bit_flash_adc clk ena rst_n ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6]
+ ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] uio_out[0] uio_out[1] uio_out[2]
+ uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] ua[0] ua[2] ua[1] VDPWR VGND uo_out[0]
.ipin clk
.ipin ena
.ipin rst_n
.ipin ua[3]
.ipin ua[4]
.ipin ua[5]
.ipin ua[6]
.ipin ua[7]
.ipin ui_in[1]
.ipin ui_in[2]
.ipin ui_in[3]
.ipin ui_in[4]
.ipin ui_in[5]
.ipin ui_in[6]
.ipin ui_in[7]
.ipin uio_in[0]
.ipin uio_in[1]
.ipin uio_in[2]
.ipin uio_in[3]
.ipin uio_in[4]
.ipin uio_in[5]
.ipin uio_in[6]
.ipin uio_in[7]
.opin uio_oe[0]
.opin uio_oe[1]
.opin uio_oe[2]
.opin uio_oe[3]
.opin uio_oe[4]
.opin uio_oe[5]
.opin uio_oe[6]
.opin uio_oe[7]
.opin uo_out[1]
.opin uo_out[2]
.opin uo_out[3]
.opin uo_out[4]
.opin uo_out[5]
.opin uo_out[6]
.opin uo_out[7]
.iopin uio_out[0]
.iopin uio_out[1]
.iopin uio_out[2]
.iopin uio_out[3]
.iopin uio_out[4]
.iopin uio_out[5]
.iopin uio_out[6]
.iopin uio_out[7]
.ipin ua[0]
.ipin ua[2]
.ipin ua[1]
.iopin VDPWR
.iopin VGND
.opin uo_out[0]
 noconn clk
 noconn ena
 noconn rst_n
 noconn ua[3]
 noconn ua[6]
 noconn #net1
 noconn ui_in[1]
 noconn ui_in[2]
 noconn ui_in[3]
 noconn ui_in[4]
 noconn ui_in[5]
 noconn ui_in[6]
 noconn ui_in[7]
 noconn uio_in[0]
 noconn uio_in[1]
 noconn uio_in[2]
 noconn uio_in[3]
 noconn uio_in[4]
 noconn uio_in[5]
 noconn uio_in[6]
 noconn uio_in[7]
 noconn uio_oe[0]
 noconn uio_oe[1]
 noconn uio_oe[2]
 noconn uio_oe[3]
 noconn uio_oe[4]
 noconn uio_oe[5]
 noconn uio_oe[6]
 noconn uio_oe[7]
 noconn uio_out[2]
 noconn uio_out[3]
 noconn uio_out[4]
 noconn uio_out[5]
 noconn uio_out[6]
 noconn uio_out[7]
 noconn ua[5]
 noconn ua[4]
 noconn ua[7]
x1 ua[0] ua[1] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] uio_out[0] uio_out[1] VDPWR VGND
+ flashADC_3bit
 noconn ua[2]
.ends

* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/adc/flashADC_3bit.sym # of pins=14
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/adc/flashADC_3bit.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/adc/flashADC_3bit.sch
.subckt flashADC_3bit vin vref dout0 dout1 dout2 d0 d1 d2 d3 d4 d5 d6 vdd vss
*.ipin vin
*.ipin vref
*.iopin vdd
*.iopin vss
*.opin dout0
*.opin dout1
*.opin dout2
*.opin d0
*.opin d1
*.opin d2
*.opin d3
*.opin d4
*.opin d5
*.opin d6
X2 vin ref0 bias_p d0 vdd vss comp_p
X3 vin ref1 bias_p d1 vdd vss comp_p
X4 vin ref2 bias_p d2 vdd vss comp_p
X5 vin ref3 bias_p d3 vdd vss comp_p
X6 vin ref4 bias_p d4 vdd vss comp_p
X7 vin ref5 bias_p d5 vdd vss comp_p
X8 vin ref6 bias_p d6 vdd vss comp_p
x9 net1 bias_p vdd vss vbias_generation
x1 d0 d1 d2 d3 d4 d5 d6 dout0 dout1 dout2 vdd vss tmux_7therm_to_3bin
x10 ref0 ref1 ref2 ref3 ref4 ref5 ref6 vref vss res_ladder_vref
* noconn #net1
.ends


* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/comparators/comp_p/comp_p.sym # of pins=6
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/comparators/comp_p/comp_p.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/comparators/comp_p/comp_p.sch
.subckt comp_p vinp vinn vbias_p vout vdd vss
*.iopin vdd
*.iopin vss
*.ipin vbias_p
*.ipin vinn
*.ipin vinp
*.opin vout
XMp_inn1 latch_left vinn tail vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XMp_inp1 latch_right vinp tail vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XMn_diode_left1 latch_left latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn_cs_left latch_right latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn_diode_right latch_right latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn_cs_right1 latch_left latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp_tail tail vbias_p vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn_out_right vout latch_right vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn_out_left out_left latch_left vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp_diode_left1 out_left out_left vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp_out vout out_left vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/vbias_generation/vbias_generation.sym # of pins=4
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/vbias_generation/vbias_generation.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/vbias_generation/vbias_generation.sch
.subckt vbias_generation bias_n bias_p vdd vss
*.opin bias_p
*.iopin vdd
*.iopin vss
*.opin bias_n
XR_bias_1 bias_1 bias_p vss sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XMn_bias bias_n bias_n vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp_bias bias_p bias_p vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR_bias_2 bias_2 bias_1 vss sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XR_bias_3 bias_3 bias_2 vss sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
XR_bias_4 bias_n bias_3 vss sky130_fd_pr__res_xhigh_po_1p41 L=7 mult=1 m=1
.ends


* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/tmux_encoder/tmux_7therm_to_3bin.sym # of pins=12
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/tmux_encoder/tmux_7therm_to_3bin.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/tmux_encoder/tmux_7therm_to_3bin.sch
.subckt tmux_7therm_to_3bin d0 d1 d2 d3 d4 d5 d6 q0 q1 q2 vdd vss
*.ipin d0
*.iopin vdd
*.opin q0
*.ipin d1
*.ipin d2
*.ipin d3
*.ipin d4
*.ipin d5
*.ipin d6
*.opin q1
*.opin q2
*.iopin vss
R1 y2 x3 sky130_fd_pr__res_generic_m1 W=1 L=1 m=1
x1 x2 x6 y2 net2 vdd vss tmux_2to1
x2 x1 x5 y2 y1 vdd vss tmux_2to1
x3 x0 x4 y2 net1 vdd vss tmux_2to1
x4 net1 net2 y1 y0 vdd vss tmux_2to1
x5 d0 x0 vdd vss buffer
x6 d1 x1 vdd vss buffer
x7 d2 x2 vdd vss buffer
x8 d3 x3 vdd vss buffer
x9 d4 x4 vdd vss buffer
x10 d5 x5 vdd vss buffer
x11 d6 x6 vdd vss buffer
x12 y0 q0 vdd vss buffer
x13 y1 q1 vdd vss buffer
x14 y2 q2 vdd vss buffer
.ends


* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/res_ladder_vref/res_ladder_vref.sym # of pins=9
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/res_ladder_vref/res_ladder_vref.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/res_ladder_vref/res_ladder_vref.sch
.subckt res_ladder_vref ref0 ref1 ref2 ref3 ref4 ref5 ref6 vref vss
*.iopin vref
*.iopin vss
*.opin ref0
*.opin ref1
*.opin ref2
*.opin ref3
*.opin ref4
*.opin ref5
*.opin ref6
XR1 ref6 vref vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR2 ref6 vref vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR3 ref5 ref6 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR4 ref4 ref5 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR5 ref3 ref4 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR6 ref2 ref3 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR7 ref1 ref2 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR8 ref0 ref1 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR9 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
XR10 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73 L=5.73 mult=1 m=1
.ends


* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/tmux/tmux_2to1.sym # of pins=6
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/tmux/tmux_2to1.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/tmux/tmux_2to1.sch
.subckt tmux_2to1 A B S Y vdd vss
*.opin Y
*.ipin S
*.iopin vss
*.iopin vdd
*.ipin A
*.ipin B
XM1 net1 S vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 net1 S vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM3 B net1 Y vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 mult=1
+ m=1
XM4 B S Y vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1 m=1
XM5 A S Y vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 mult=1
+ m=1
XM6 A net1 Y vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
.ends


* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/buffer/buffer.sym # of pins=4
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/buffer/buffer.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/buffer/buffer.sch
.subckt buffer in out vdd vss
*.ipin in
*.opin out
*.iopin vdd
*.iopin vss
X1 in net1 vdd vss inv
X2 net1 out vdd vss inv
.ends


* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/inv/inv.sym # of pins=4
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/inv/inv.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/inv/inv.sch
.subckt inv vin vout vdd vss
*.ipin vin
*.opin vout
*.ipin vdd
*.ipin vss
XMn vout vin vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XMp vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends

.end
