** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/buffer/buffer.sch
.subckt buffer vdd in out vss
*.ipin in
*.opin out
*.iopin vdd
*.iopin vss
X1 in net1 vdd vss inv
X2 net1 out vdd vss inv
**.ends

* expanding   symbol:  /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/inv/inv.sym # of pins=4
** sym_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/inv/inv.sym
** sch_path: /home/bmott/ttsky25b_tiny_chaos/xsch/ip/logic/inv/inv.sch
.subckt inv vin vout vdd vss
*.ipin vin
*.opin vout
*.ipin vdd
*.ipin vss
XMn vout vin vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XMp vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends

.end
