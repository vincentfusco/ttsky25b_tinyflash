magic
tech sky130A
magscale 1 2
timestamp 1762640459
<< nwell >>
rect 1854 622 2908 1460
rect 1854 -2294 2908 -1456
rect 3060 -1502 3510 -1394
rect 800 -5210 3750 -3534
rect 800 -8126 3750 -6450
<< pwell >>
rect 1770 -104 2908 622
rect 800 -2864 3750 -2294
rect 800 -2972 3056 -2864
rect 3506 -2972 3750 -2864
rect 800 -3534 3750 -2972
rect 800 -6450 3750 -5210
rect 800 -8746 3750 -8126
<< metal1 >>
rect -42 1448 3750 1460
rect -42 1394 -26 1448
rect 3720 1394 3750 1448
rect -42 1380 3750 1394
rect -42 582 198 662
rect 3648 582 3740 662
rect -42 60 3750 82
rect -42 -44 -18 60
rect 3720 -44 3750 60
rect -42 -48 248 -44
rect 698 -48 3750 -44
rect -42 -78 3750 -48
rect -42 -658 198 -578
rect 1038 -782 1040 -466
rect 3648 -658 3740 -578
rect -42 -1398 3750 -1376
rect -42 -1502 -18 -1398
rect 3720 -1502 3750 -1398
rect -42 -1536 3750 -1502
rect -42 -2334 198 -2254
rect 2666 -2254 2802 -2238
rect 2666 -2262 2972 -2254
rect 2666 -2406 2684 -2262
rect 2790 -2334 2972 -2262
rect 3648 -2334 3740 -2254
rect 2790 -2406 2802 -2334
rect 2666 -2426 2802 -2406
rect -42 -2858 3750 -2834
rect -42 -2864 244 -2858
rect 694 -2864 3750 -2858
rect -42 -2968 -20 -2864
rect 3718 -2968 3750 -2864
rect -42 -2994 3750 -2968
rect 916 -3074 1116 -3044
rect 916 -3184 942 -3074
rect 1082 -3184 1116 -3074
rect 916 -3216 1116 -3184
rect 916 -3494 1116 -3450
rect -42 -3574 198 -3494
rect 698 -3574 1116 -3494
rect -42 -4318 3750 -4292
rect -42 -4422 -22 -4318
rect 3716 -4422 3750 -4318
rect -42 -4452 3750 -4422
rect -42 -5250 198 -5170
rect -42 -5774 3750 -5750
rect -42 -5776 242 -5774
rect 692 -5776 3750 -5774
rect -42 -5880 -24 -5776
rect 3714 -5880 3750 -5776
rect -42 -5882 242 -5880
rect 692 -5882 3750 -5880
rect -42 -5910 3750 -5882
rect -42 -6490 198 -6410
rect -42 -7238 3750 -7208
rect -42 -7342 -22 -7238
rect 3716 -7342 3750 -7238
rect -42 -7368 3750 -7342
rect -42 -8166 198 -8086
rect -42 -8678 3750 -8666
rect -42 -8732 -26 -8678
rect 3720 -8732 3750 -8678
rect -42 -8738 232 -8732
rect 722 -8738 3750 -8732
rect -42 -8746 3750 -8738
<< via1 >>
rect -26 1394 3720 1448
rect 640 872 704 1200
rect 1216 882 1280 1210
rect 1702 958 1760 1190
rect 1446 776 1524 878
rect 982 456 1038 624
rect 2968 596 3124 648
rect -18 -44 3720 60
rect 248 -48 698 -44
rect 2264 -374 2322 -244
rect 980 -782 1038 -466
rect 2506 -480 2572 -252
rect 2758 -372 2816 -242
rect 2036 -740 2092 -490
rect 2968 -644 3126 -590
rect 642 -1196 706 -868
rect 1216 -1202 1280 -874
rect 1446 -900 1524 -754
rect 1696 -1162 1766 -906
rect -18 -1502 3720 -1398
rect 644 -2040 712 -1930
rect 1212 -2044 1276 -1896
rect 1434 -1900 1528 -1734
rect 1698 -2040 1760 -1912
rect 984 -2450 1038 -2134
rect 2684 -2406 2790 -2262
rect 244 -2864 694 -2858
rect -20 -2968 3718 -2864
rect 942 -3184 1082 -3074
rect -22 -4422 3716 -4318
rect 646 -4942 704 -4656
rect 242 -5776 692 -5774
rect -24 -5880 3714 -5776
rect 242 -5882 692 -5880
rect 642 -7010 708 -6726
rect -22 -7342 3716 -7238
rect 642 -7858 704 -7578
rect -26 -8732 3720 -8678
rect 232 -8738 722 -8732
<< metal2 >>
rect -42 1450 3750 1460
rect -42 1448 226 1450
rect 716 1448 3750 1450
rect -42 1394 -26 1448
rect 3720 1394 3750 1448
rect -42 1390 226 1394
rect 716 1390 3750 1394
rect -42 1380 3750 1390
rect 1208 1210 1288 1218
rect 628 1200 714 1210
rect 628 872 640 1200
rect 704 1018 714 1200
rect 1208 1018 1216 1210
rect 704 946 1216 1018
rect 704 872 714 946
rect 1208 882 1216 946
rect 1280 882 1288 1210
rect 1692 1190 1770 1200
rect 1692 958 1702 1190
rect 1760 958 1770 1190
rect 1692 948 1770 958
rect 1208 872 1288 882
rect 1428 888 2334 892
rect 1428 878 2264 888
rect 628 860 714 872
rect 1428 776 1446 878
rect 1524 816 2264 878
rect 2324 816 2334 888
rect 1524 812 2334 816
rect 1524 776 1542 812
rect 1428 760 1542 776
rect 2496 654 3132 664
rect 978 624 1044 634
rect 978 456 982 624
rect 1038 456 1044 624
rect 2496 598 2502 654
rect 2576 648 3132 654
rect 2576 598 2968 648
rect 2496 596 2968 598
rect 3124 596 3132 648
rect 2496 588 3132 596
rect 978 446 1044 456
rect -42 60 3750 82
rect -42 -44 -18 60
rect 3720 -44 3750 60
rect -42 -48 248 -44
rect 698 -48 3048 -44
rect 3498 -48 3750 -44
rect -42 -78 3750 -48
rect 2254 -244 2334 -238
rect 2254 -374 2264 -244
rect 2322 -374 2334 -244
rect 2254 -378 2334 -374
rect 2496 -252 2584 -240
rect 980 -460 1042 -456
rect 970 -466 1050 -460
rect 970 -782 980 -466
rect 1038 -782 1050 -466
rect 2032 -490 2098 -442
rect 2496 -480 2506 -252
rect 2572 -480 2584 -252
rect 2748 -242 2826 -232
rect 2748 -372 2758 -242
rect 2816 -372 2826 -242
rect 2748 -382 2826 -372
rect 2496 -490 2584 -480
rect 2032 -740 2036 -490
rect 2092 -740 2098 -490
rect 2032 -746 2098 -740
rect 2948 -590 3148 -578
rect 2948 -644 2968 -590
rect 3126 -644 3148 -590
rect 2948 -658 3148 -644
rect 2948 -746 3004 -658
rect 970 -794 1050 -782
rect 1438 -754 3004 -746
rect 630 -868 716 -858
rect 630 -1196 642 -868
rect 706 -984 716 -868
rect 1204 -874 1290 -862
rect 1204 -984 1216 -874
rect 706 -1064 1216 -984
rect 706 -1196 716 -1064
rect 630 -1206 716 -1196
rect 1204 -1202 1216 -1064
rect 1280 -1202 1290 -874
rect 1438 -900 1446 -754
rect 1524 -812 3004 -754
rect 1524 -900 1532 -812
rect 1438 -908 1532 -900
rect 1686 -906 1776 -888
rect 1686 -1162 1696 -906
rect 1766 -1162 1776 -906
rect 1686 -1174 1776 -1162
rect 1204 -1210 1290 -1202
rect -42 -1398 3750 -1376
rect -42 -1502 -18 -1398
rect 3720 -1502 3750 -1398
rect -42 -1514 246 -1502
rect 696 -1514 3750 -1502
rect -42 -1536 3750 -1514
rect 1424 -1724 2824 -1714
rect 1424 -1734 2756 -1724
rect 1206 -1896 1284 -1886
rect 634 -1930 722 -1914
rect 634 -2040 644 -1930
rect 712 -1984 722 -1930
rect 1206 -1984 1212 -1896
rect 712 -2040 1212 -1984
rect 634 -2044 1212 -2040
rect 1276 -2044 1284 -1896
rect 1424 -1900 1434 -1734
rect 1528 -1804 2756 -1734
rect 2816 -1804 2824 -1724
rect 1528 -1814 2824 -1804
rect 1528 -1900 1540 -1814
rect 1424 -1918 1540 -1900
rect 1686 -1912 1772 -1902
rect 634 -2054 1284 -2044
rect 1686 -2040 1698 -1912
rect 1760 -2040 1772 -1912
rect 1686 -2052 1772 -2040
rect 978 -2134 1044 -2118
rect 978 -2450 982 -2134
rect 1038 -2450 1044 -2134
rect 978 -2538 1044 -2450
rect 2666 -2262 2802 -2236
rect 2666 -2406 2684 -2262
rect 2790 -2406 2802 -2262
rect 2666 -2426 2802 -2406
rect 2666 -2538 2732 -2426
rect 978 -2606 2732 -2538
rect -42 -2858 3750 -2834
rect -42 -2864 244 -2858
rect 694 -2864 3052 -2858
rect 3516 -2864 3750 -2858
rect -42 -2968 -20 -2864
rect 3718 -2968 3750 -2864
rect -42 -2994 3750 -2968
rect 922 -3074 1100 -3062
rect 922 -3184 942 -3074
rect 1082 -3184 1100 -3074
rect 922 -3196 1100 -3184
rect -42 -4312 3750 -4292
rect -42 -4318 254 -4312
rect 704 -4318 3750 -4312
rect -42 -4422 -22 -4318
rect 3716 -4422 3750 -4318
rect -42 -4452 3750 -4422
rect 634 -4656 716 -4640
rect 634 -4942 646 -4656
rect 704 -4748 716 -4656
rect 1536 -4644 1614 -4628
rect 1536 -4748 1550 -4644
rect 704 -4820 1550 -4748
rect 1606 -4820 1614 -4644
rect 704 -4830 1614 -4820
rect 704 -4942 716 -4830
rect 634 -4954 716 -4942
rect -42 -5774 3750 -5750
rect -42 -5776 242 -5774
rect 692 -5776 3038 -5774
rect 3502 -5776 3750 -5774
rect -42 -5880 -24 -5776
rect 3714 -5880 3750 -5776
rect -42 -5882 242 -5880
rect 692 -5882 3038 -5880
rect 3502 -5882 3750 -5880
rect -42 -5910 3750 -5882
rect 630 -6726 720 -6710
rect 630 -7010 642 -6726
rect 708 -6830 720 -6726
rect 708 -6842 1452 -6830
rect 708 -6904 1216 -6842
rect 1444 -6904 1452 -6842
rect 708 -6914 1452 -6904
rect 708 -7010 720 -6914
rect 630 -7024 720 -7010
rect -42 -7234 3750 -7208
rect -42 -7238 242 -7234
rect 692 -7238 3750 -7234
rect -42 -7342 -22 -7238
rect 3716 -7342 3750 -7238
rect -42 -7368 3750 -7342
rect 628 -7578 714 -7564
rect 628 -7858 642 -7578
rect 704 -7786 714 -7578
rect 704 -7796 1766 -7786
rect 704 -7858 1482 -7796
rect 628 -7866 1482 -7858
rect 1756 -7866 1766 -7796
rect 628 -7874 1766 -7866
rect -42 -8676 3750 -8666
rect -42 -8678 3032 -8676
rect 3522 -8678 3750 -8676
rect -42 -8732 -26 -8678
rect 3720 -8732 3750 -8678
rect -42 -8738 232 -8732
rect 722 -8736 3032 -8732
rect 3522 -8736 3750 -8732
rect 722 -8738 3750 -8736
rect -42 -8746 3750 -8738
<< via2 >>
rect 226 1448 716 1450
rect 226 1394 716 1448
rect 226 1390 716 1394
rect 1702 958 1760 1190
rect 2264 816 2324 888
rect 982 456 1038 624
rect 2502 598 2576 654
rect 3048 -44 3498 60
rect 3048 -48 3498 -44
rect 2264 -374 2322 -244
rect 980 -782 1038 -466
rect 2506 -478 2572 -252
rect 2758 -372 2816 -242
rect 1696 -1162 1766 -906
rect 246 -1502 696 -1406
rect 2124 -1500 2538 -1404
rect 246 -1514 696 -1502
rect 2756 -1804 2816 -1724
rect 1698 -2040 1760 -1912
rect 982 -2450 984 -2134
rect 984 -2450 1038 -2134
rect 3052 -2864 3516 -2858
rect 3052 -2966 3516 -2864
rect 942 -3184 1082 -3074
rect 254 -4318 704 -4312
rect 254 -4420 704 -4318
rect 2130 -4418 2544 -4322
rect 1550 -4820 1606 -4644
rect 3038 -5776 3502 -5774
rect 3038 -5880 3502 -5776
rect 3038 -5882 3502 -5880
rect 1216 -6904 1444 -6842
rect 242 -7238 692 -7234
rect 242 -7342 692 -7238
rect 2118 -7342 2532 -7246
rect 1482 -7866 1756 -7796
rect 3032 -8678 3522 -8676
rect 3032 -8732 3522 -8678
rect 3032 -8736 3522 -8732
<< metal3 >>
rect 218 1450 738 1460
rect 218 1390 226 1450
rect 716 1390 738 1450
rect 218 -1406 738 1390
rect 1692 1190 1770 1200
rect 1692 958 1702 1190
rect 1760 1004 1770 1190
rect 1760 958 1942 1004
rect 1692 906 1942 958
rect 218 -1514 246 -1406
rect 696 -1514 738 -1406
rect 218 -4312 738 -1514
rect 974 624 1044 634
rect 974 456 982 624
rect 1038 456 1044 624
rect 974 -466 1044 456
rect 974 -782 980 -466
rect 1038 -782 1044 -466
rect 974 -2134 1044 -782
rect 1686 -906 1772 -898
rect 974 -2450 982 -2134
rect 1038 -2450 1044 -2134
rect 974 -3064 1044 -2450
rect 1376 -1090 1452 -1088
rect 1686 -1090 1696 -906
rect 1376 -1162 1696 -1090
rect 1766 -1162 1772 -906
rect 1376 -1174 1772 -1162
rect 932 -3074 1092 -3064
rect 932 -3184 942 -3074
rect 1082 -3184 1092 -3074
rect 932 -3190 1092 -3184
rect 218 -4420 254 -4312
rect 704 -4420 738 -4312
rect 218 -7234 738 -4420
rect 1376 -6830 1452 -1174
rect 1864 -1316 1942 906
rect 2258 888 2334 898
rect 2258 816 2264 888
rect 2324 816 2334 888
rect 2258 -244 2334 816
rect 2258 -374 2264 -244
rect 2322 -374 2334 -244
rect 2258 -382 2334 -374
rect 2496 654 2584 664
rect 2496 598 2502 654
rect 2576 598 2584 654
rect 2496 -252 2584 598
rect 3016 60 3564 1460
rect 3016 -48 3048 60
rect 3498 -48 3564 60
rect 2496 -478 2506 -252
rect 2572 -478 2584 -252
rect 2496 -488 2584 -478
rect 2750 -242 2824 -234
rect 2750 -372 2758 -242
rect 2816 -372 2824 -242
rect 1536 -1380 1942 -1316
rect 1536 -4644 1614 -1380
rect 2032 -1404 2622 -1376
rect 2032 -1500 2124 -1404
rect 2538 -1500 2622 -1404
rect 1536 -4820 1550 -4644
rect 1606 -4820 1614 -4644
rect 1536 -4830 1614 -4820
rect 1692 -1912 1766 -1906
rect 1692 -2040 1698 -1912
rect 1760 -2040 1766 -1912
rect 1194 -6842 1452 -6830
rect 1194 -6904 1216 -6842
rect 1444 -6904 1452 -6842
rect 1194 -6914 1452 -6904
rect 218 -7342 242 -7234
rect 692 -7342 738 -7234
rect 218 -8746 738 -7342
rect 1692 -7786 1766 -2040
rect 1466 -7796 1766 -7786
rect 1466 -7866 1482 -7796
rect 1756 -7866 1766 -7796
rect 1466 -7874 1766 -7866
rect 2032 -4322 2622 -1500
rect 2750 -1724 2824 -372
rect 2750 -1804 2756 -1724
rect 2816 -1804 2824 -1724
rect 2750 -1814 2824 -1804
rect 2032 -4418 2130 -4322
rect 2544 -4418 2622 -4322
rect 2032 -7246 2622 -4418
rect 2032 -7342 2118 -7246
rect 2532 -7342 2622 -7246
rect 2032 -8746 2622 -7342
rect 3016 -2858 3564 -48
rect 3016 -2966 3052 -2858
rect 3516 -2966 3564 -2858
rect 3016 -5774 3564 -2966
rect 3016 -5882 3038 -5774
rect 3502 -5882 3564 -5774
rect 3016 -8676 3564 -5882
rect 3016 -8736 3032 -8676
rect 3522 -8736 3564 -8676
rect 3016 -8746 3564 -8736
use buffer  buffer_0
timestamp 1762640459
transform 1 0 178 0 1 -18
box -220 20 622 1478
use buffer  buffer_1
timestamp 1762640459
transform 1 0 178 0 -1 22
box -220 20 622 1478
use buffer  buffer_2
timestamp 1762640459
transform 1 0 178 0 1 -2934
box -220 20 622 1478
use buffer  buffer_3
timestamp 1762640459
transform 1 0 178 0 -1 -2894
box -220 20 622 1478
use buffer  buffer_4
timestamp 1762640459
transform 1 0 178 0 1 -5850
box -220 20 622 1478
use buffer  buffer_5
timestamp 1762640459
transform 1 0 178 0 -1 -5810
box -220 20 622 1478
use buffer  buffer_6
timestamp 1762640459
transform 1 0 178 0 1 -8766
box -220 20 622 1478
use buffer  buffer_7
timestamp 1762640459
transform 1 0 3128 0 1 -18
box -220 20 622 1478
use buffer  buffer_8
timestamp 1762640459
transform 1 0 3128 0 -1 22
box -220 20 622 1478
use buffer  buffer_9
timestamp 1762640459
transform 1 0 3128 0 1 -2934
box -220 20 622 1478
use sky130_fd_pr__res_generic_m1_SPQYYJ  R1
timestamp 1762640459
transform 1 0 1016 0 1 -3335
box -100 -157 100 157
use tmux_2to1  tmux_2to1_0
timestamp 1762640459
transform 1 0 714 0 1 588
box 86 -586 1140 872
use tmux_2to1  tmux_2to1_1
timestamp 1762640459
transform 1 0 714 0 -1 -584
box 86 -586 1140 872
use tmux_2to1  tmux_2to1_2
timestamp 1762640459
transform 1 0 714 0 1 -2328
box 86 -586 1140 872
use tmux_2to1  tmux_2to1_3
timestamp 1762640459
transform 1 0 1768 0 -1 -584
box 86 -586 1140 872
<< labels >>
rlabel metal1 -42 582 198 662 1 d0
port 0 n
rlabel metal1 -42 -658 198 -578 1 d1
port 1 n
rlabel metal1 -42 -2334 198 -2254 1 d2
port 2 n
rlabel metal1 -42 -3574 198 -3494 1 d3
port 3 n
rlabel metal1 -42 -5250 198 -5170 1 d4
port 4 n
rlabel metal1 -42 -6490 198 -6410 1 d5
port 5 n
rlabel metal1 -42 -8166 198 -8086 1 d6
port 6 n
rlabel metal1 3648 582 3740 662 1 q0
port 7 n
rlabel metal1 3648 -658 3740 -578 1 q1
port 8 n
rlabel metal1 3648 -2334 3740 -2254 1 q2
port 9 n
rlabel metal3 218 -1406 738 1390 1 vdd
port 10 n
rlabel metal3 3016 60 3536 1460 1 vss
port 11 n
<< end >>
