* NGSPICE file created from tmux_7therm_to_3bin_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_A6MZLZ B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 S B 0.14266f
C1 D G 0.02934f
C2 S D 0.32105f
C3 D B 0.14266f
C4 S G 0.02934f
C5 B G 0.24043f
C6 S VSUBS 0.09023f
C7 D VSUBS 0.09023f
C8 G VSUBS 0.11914f
C9 B VSUBS 1.5811f
.ends

.subckt sky130_fd_pr__nfet_01v8_MH3LLV B D S G
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 S D 0.16211f
C1 S G 0.02545f
C2 G D 0.02545f
C3 S B 0.1317f
C4 D B 0.1317f
C5 G B 0.34289f
.ends

.subckt tmux_2to1 Y vdd XM5/G B A S vss
XXM1 vdd vdd XM5/G S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM2 vss vss XM5/G S sky130_fd_pr__nfet_01v8_MH3LLV
XXM3 vdd A Y S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM4 vss A Y XM5/G sky130_fd_pr__nfet_01v8_MH3LLV
XXM5 vdd Y B XM5/G vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM6 vss Y B S sky130_fd_pr__nfet_01v8_MH3LLV
C0 vdd Y 0.18933f
C1 vdd XM5/G 0.17343f
C2 vdd A 0.05809f
C3 B Y 0.03022f
C4 S Y 0.13093f
C5 B XM5/G 0.09611f
C6 S XM5/G 0.4752f
C7 S A 0.09932f
C8 XM5/G Y 0.31571f
C9 A Y 0.03022f
C10 XM5/G A 0.66126f
C11 B vdd 0.11322f
C12 vdd S 0.27839f
C13 B S 0.0426f
C14 B vss 0.39578f
C15 S vss 1.22376f
C16 Y vss 0.38976f
C17 XM5/G vss 0.68597f
C18 vdd vss 4.09633f
C19 A vss 0.18036f
.ends

.subckt sky130_fd_pr__res_generic_m1_SPQYYJ R1 R2 m1_n100_n100# VSUBS
R0 R1 R2 sky130_fd_pr__res_generic_m1 w=1 l=1
C0 R2 VSUBS 0.07104f
C1 R1 VSUBS 0.07104f
C2 m1_n100_n100# VSUBS 0.10692f
.ends

.subckt inv vin vdd vout vss
XXMn vss vss vout vin sky130_fd_pr__nfet_01v8_MH3LLV
XXMp vdd vdd vout vin vss sky130_fd_pr__pfet_01v8_A6MZLZ
C0 vdd vin 0.13776f
C1 vdd vout 0.11998f
C2 vout vin 0.12658f
C3 vin vss 0.56678f
C4 vout vss 0.40687f
C5 vdd vss 1.84972f
.ends

.subckt buffer in out vdd inv_1/vin vss
Xinv_0 in vdd inv_1/vin vss inv
Xinv_1 inv_1/vin vdd out vss inv
C0 vdd in 0.01965f
C1 out inv_1/vin 0.0071f
C2 vdd inv_1/vin 0.16476f
C3 in inv_1/vin 0.01628f
C4 vdd out 0.00589f
C5 inv_1/vin vss 0.60193f
C6 out vss 0.3255f
C7 in vss 0.41789f
C8 vdd vss 3.06334f
.ends

.subckt tmux_7therm_to_3bin_extracted d0 d1 d2 d3 d4 d5 d6 q0 q1 q2 vdd vss
Xtmux_2to1_1 buffer_8/in vdd tmux_2to1_1/XM5/G buffer_5/out buffer_1/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_2 tmux_2to1_3/B vdd tmux_2to1_2/XM5/G buffer_6/out buffer_2/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_3 buffer_7/in vdd tmux_2to1_3/XM5/G tmux_2to1_3/B tmux_2to1_3/A buffer_8/in
+ vss tmux_2to1
XR1 R1/R1 R1/R2 R1/m1_n100_n100# vss sky130_fd_pr__res_generic_m1_SPQYYJ
Xbuffer_0 d0 buffer_0/out vdd buffer_0/inv_1/vin vss buffer
Xbuffer_1 d1 buffer_1/out vdd buffer_1/inv_1/vin vss buffer
Xbuffer_2 d2 buffer_2/out vdd buffer_2/inv_1/vin vss buffer
Xbuffer_3 d3 R1/R2 vdd buffer_3/inv_1/vin vss buffer
Xbuffer_4 d4 buffer_4/out vdd buffer_4/inv_1/vin vss buffer
Xbuffer_5 d5 buffer_5/out vdd buffer_5/inv_1/vin vss buffer
Xbuffer_6 d6 buffer_6/out vdd buffer_6/inv_1/vin vss buffer
Xbuffer_7 buffer_7/in q0 vdd buffer_7/inv_1/vin vss buffer
Xbuffer_8 buffer_8/in q1 vdd buffer_8/inv_1/vin vss buffer
Xbuffer_9 R1/R1 q2 vdd buffer_9/inv_1/vin vss buffer
Xtmux_2to1_0 tmux_2to1_3/A vdd tmux_2to1_0/XM5/G buffer_4/out buffer_0/out R1/R1 vss
+ tmux_2to1
X0 buffer_4/inv_1/vin d4.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X1 buffer_1/inv_1/vin d1.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X2 buffer_1/inv_1/vin d1.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X3 buffer_5/inv_1/vin d5.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X4 buffer_3/inv_1/vin d3.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X5 buffer_5/inv_1/vin d5.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X6 buffer_0/inv_1/vin d0.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X7 buffer_3/inv_1/vin d3.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X8 buffer_4/inv_1/vin d4.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X9 buffer_2/inv_1/vin d2.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X10 buffer_0/inv_1/vin d0.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X11 buffer_6/inv_1/vin d6.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X12 buffer_2/inv_1/vin d2.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X13 buffer_6/inv_1/vin d6.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
R0 vdd.n71 vdd.n59 1789.41
R1 vdd.n68 vdd.n59 1789.41
R2 vdd.n71 vdd.n60 1789.41
R3 vdd.n77 vdd.n54 1789.41
R4 vdd.n74 vdd.n54 1789.41
R5 vdd.n77 vdd.n55 1789.41
R6 vdd.n74 vdd.n55 1789.41
R7 vdd.n41 vdd.n12 1789.41
R8 vdd.n41 vdd.n13 1789.41
R9 vdd.n81 vdd.n5 1789.41
R10 vdd.n52 vdd.n5 1789.41
R11 vdd.n34 vdd.n15 1789.41
R12 vdd.n37 vdd.n15 1789.41
R13 vdd.n34 vdd.n16 1789.41
R14 vdd.n37 vdd.n16 1789.41
R15 vdd.n31 vdd.n20 1789.41
R16 vdd.n28 vdd.n21 1789.41
R17 vdd.n31 vdd.n21 1789.41
R18 vdd.n124 vdd.n98 1789.41
R19 vdd.n98 vdd.n94 1789.41
R20 vdd.n124 vdd.n99 1789.41
R21 vdd.n99 vdd.n94 1789.41
R22 vdd.n97 vdd.n91 1789.41
R23 vdd.n126 vdd.n91 1789.41
R24 vdd.n97 vdd.n92 1789.41
R25 vdd.n126 vdd.n92 1789.41
R26 vdd.n107 vdd.n102 1789.41
R27 vdd.n116 vdd.n102 1789.41
R28 vdd.n107 vdd.n103 1789.41
R29 vdd.n116 vdd.n103 1789.41
R30 vdd.n109 vdd.n105 1789.41
R31 vdd.n114 vdd.n109 1789.41
R32 vdd.n110 vdd.n105 1789.41
R33 vdd.n114 vdd.n110 1789.41
R34 vdd.n208 vdd.n193 1789.41
R35 vdd.n215 vdd.n193 1789.41
R36 vdd.n208 vdd.n194 1789.41
R37 vdd.n215 vdd.n194 1789.41
R38 vdd.n224 vdd.n186 1789.41
R39 vdd.n205 vdd.n186 1789.41
R40 vdd.n224 vdd.n187 1789.41
R41 vdd.n205 vdd.n187 1789.41
R42 vdd.n336 vdd.n329 1789.41
R43 vdd.n329 vdd.n327 1789.41
R44 vdd.n348 vdd.n181 1789.41
R45 vdd.n350 vdd.n181 1789.41
R46 vdd.n310 vdd.n291 1789.41
R47 vdd.n310 vdd.n292 1789.41
R48 vdd.n324 vdd.n250 1789.41
R49 vdd.n324 vdd.n251 1789.41
R50 vdd.n284 vdd.n256 1789.41
R51 vdd.n313 vdd.n256 1789.41
R52 vdd.n284 vdd.n257 1789.41
R53 vdd.n313 vdd.n257 1789.41
R54 vdd.n276 vdd.n268 1789.41
R55 vdd.n268 vdd.n263 1789.41
R56 vdd.n276 vdd.n269 1789.41
R57 vdd.n269 vdd.n263 1789.41
R58 vdd.n210 vdd.n196 1789.41
R59 vdd.n213 vdd.n196 1789.41
R60 vdd.n210 vdd.n197 1789.41
R61 vdd.n213 vdd.n197 1789.41
R62 vdd.n199 vdd.n184 1789.41
R63 vdd.n204 vdd.n199 1789.41
R64 vdd.n200 vdd.n184 1789.41
R65 vdd.n204 vdd.n200 1789.41
R66 vdd.n328 vdd.n247 1789.41
R67 vdd.n338 vdd.n247 1789.41
R68 vdd.n243 vdd.n227 1789.41
R69 vdd.n243 vdd.n183 1789.41
R70 vdd.n286 vdd.n259 1789.41
R71 vdd.n289 vdd.n259 1789.41
R72 vdd.n286 vdd.n260 1789.41
R73 vdd.n289 vdd.n260 1789.41
R74 vdd.n278 vdd.n264 1789.41
R75 vdd.n281 vdd.n264 1789.41
R76 vdd.n278 vdd.n265 1789.41
R77 vdd.n281 vdd.n265 1789.41
R78 vdd.n167 vdd.n141 1789.41
R79 vdd.n141 vdd.n137 1789.41
R80 vdd.n167 vdd.n142 1789.41
R81 vdd.n142 vdd.n137 1789.41
R82 vdd.n140 vdd.n134 1789.41
R83 vdd.n169 vdd.n134 1789.41
R84 vdd.n140 vdd.n135 1789.41
R85 vdd.n169 vdd.n135 1789.41
R86 vdd.n150 vdd.n145 1789.41
R87 vdd.n159 vdd.n145 1789.41
R88 vdd.n150 vdd.n146 1789.41
R89 vdd.n159 vdd.n146 1789.41
R90 vdd.n152 vdd.n148 1789.41
R91 vdd.n157 vdd.n152 1789.41
R92 vdd.n153 vdd.n148 1789.41
R93 vdd.n157 vdd.n153 1789.41
R94 vdd.n40 vdd.n38 1315.04
R95 vdd.n7 vdd.n4 1231.76
R96 vdd.n8 vdd.n7 1231.76
R97 vdd.n47 vdd.n46 1231.76
R98 vdd.n46 vdd.n10 1231.76
R99 vdd.n229 vdd.n228 1231.76
R100 vdd.n228 vdd.n180 1231.76
R101 vdd.n331 vdd.n231 1231.76
R102 vdd.n331 vdd.n330 1231.76
R103 vdd.n300 vdd.n299 1231.76
R104 vdd.n299 vdd.n298 1231.76
R105 vdd.n305 vdd.n294 1231.76
R106 vdd.n305 vdd.n295 1231.76
R107 vdd.n239 vdd.n236 1231.76
R108 vdd.n239 vdd.n238 1231.76
R109 vdd.n340 vdd.n235 1231.76
R110 vdd.n340 vdd.n339 1231.76
R111 vdd.n47 vdd.n12 557.648
R112 vdd.n48 vdd.n47 557.648
R113 vdd.n48 vdd.n4 557.648
R114 vdd.n81 vdd.n4 557.648
R115 vdd.n13 vdd.n10 557.648
R116 vdd.n50 vdd.n10 557.648
R117 vdd.n50 vdd.n8 557.648
R118 vdd.n52 vdd.n8 557.648
R119 vdd.n336 vdd.n231 557.648
R120 vdd.n346 vdd.n231 557.648
R121 vdd.n346 vdd.n229 557.648
R122 vdd.n348 vdd.n229 557.648
R123 vdd.n330 vdd.n327 557.648
R124 vdd.n330 vdd.n233 557.648
R125 vdd.n233 vdd.n180 557.648
R126 vdd.n350 vdd.n180 557.648
R127 vdd.n294 vdd.n291 557.648
R128 vdd.n302 vdd.n294 557.648
R129 vdd.n302 vdd.n300 557.648
R130 vdd.n300 vdd.n250 557.648
R131 vdd.n295 vdd.n292 557.648
R132 vdd.n296 vdd.n295 557.648
R133 vdd.n298 vdd.n296 557.648
R134 vdd.n298 vdd.n251 557.648
R135 vdd.n328 vdd.n235 557.648
R136 vdd.n344 vdd.n235 557.648
R137 vdd.n344 vdd.n236 557.648
R138 vdd.n236 vdd.n227 557.648
R139 vdd.n339 vdd.n338 557.648
R140 vdd.n339 vdd.n234 557.648
R141 vdd.n238 vdd.n234 557.648
R142 vdd.n238 vdd.n183 557.648
R143 vdd.n70 vdd.n61 190.871
R144 vdd.n70 vdd 190.871
R145 vdd vdd.n69 190.871
R146 vdd.n76 vdd.n56 190.871
R147 vdd.n76 vdd 190.871
R148 vdd vdd.n75 190.871
R149 vdd.n43 vdd.n42 190.871
R150 vdd.n42 vdd 190.871
R151 vdd.n82 vdd.n3 190.871
R152 vdd vdd.n3 190.871
R153 vdd.n35 vdd.n18 190.871
R154 vdd vdd.n35 190.871
R155 vdd.n36 vdd 190.871
R156 vdd.n30 vdd 190.871
R157 vdd vdd.n29 190.871
R158 vdd.n29 vdd.n26 190.871
R159 vdd.n123 vdd 190.871
R160 vdd.n100 vdd 190.871
R161 vdd.n123 vdd.n122 190.871
R162 vdd.n96 vdd 190.871
R163 vdd.n127 vdd 190.871
R164 vdd.n96 vdd.n90 190.871
R165 vdd.n106 vdd.n101 190.871
R166 vdd.n106 vdd 190.871
R167 vdd.n117 vdd 190.871
R168 vdd.n113 vdd 190.871
R169 vdd vdd.n112 190.871
R170 vdd.n112 vdd.n111 190.871
R171 vdd.n207 vdd 190.871
R172 vdd.n216 vdd 190.871
R173 vdd.n207 vdd.n192 190.871
R174 vdd.n223 vdd 190.871
R175 vdd.n188 vdd 190.871
R176 vdd.n223 vdd.n222 190.871
R177 vdd vdd.n335 190.871
R178 vdd.n335 vdd.n334 190.871
R179 vdd vdd.n179 190.871
R180 vdd.n351 vdd.n179 190.871
R181 vdd.n309 vdd 190.871
R182 vdd.n309 vdd.n308 190.871
R183 vdd.n323 vdd 190.871
R184 vdd.n323 vdd.n322 190.871
R185 vdd.n283 vdd 190.871
R186 vdd.n314 vdd 190.871
R187 vdd.n283 vdd.n255 190.871
R188 vdd.n275 vdd 190.871
R189 vdd.n270 vdd 190.871
R190 vdd.n275 vdd.n274 190.871
R191 vdd.n211 vdd.n198 190.871
R192 vdd vdd.n211 190.871
R193 vdd.n212 vdd 190.871
R194 vdd.n202 vdd.n201 190.871
R195 vdd vdd.n202 190.871
R196 vdd.n203 vdd 190.871
R197 vdd.n248 vdd.n237 190.871
R198 vdd vdd.n248 190.871
R199 vdd.n244 vdd.n242 190.871
R200 vdd vdd.n244 190.871
R201 vdd.n287 vdd.n261 190.871
R202 vdd vdd.n287 190.871
R203 vdd.n288 vdd 190.871
R204 vdd.n280 vdd 190.871
R205 vdd vdd.n279 190.871
R206 vdd.n279 vdd.n267 190.871
R207 vdd.n166 vdd 190.871
R208 vdd.n143 vdd 190.871
R209 vdd.n166 vdd.n165 190.871
R210 vdd.n139 vdd 190.871
R211 vdd.n170 vdd 190.871
R212 vdd.n139 vdd.n133 190.871
R213 vdd.n149 vdd.n144 190.871
R214 vdd.n149 vdd 190.871
R215 vdd.n160 vdd 190.871
R216 vdd.n156 vdd 190.871
R217 vdd vdd.n155 190.871
R218 vdd.n155 vdd.n154 190.871
R219 vdd.n69 vdd.n66 190.494
R220 vdd.n75 vdd.n57 190.494
R221 vdd.n36 vdd.n17 190.494
R222 vdd.n30 vdd.n25 190.494
R223 vdd.n121 vdd.n100 190.494
R224 vdd.n128 vdd.n127 190.494
R225 vdd.n118 vdd.n117 190.494
R226 vdd.n113 vdd.n88 190.494
R227 vdd.n217 vdd.n216 190.494
R228 vdd.n221 vdd.n188 190.494
R229 vdd.n315 vdd.n314 190.494
R230 vdd.n273 vdd.n270 190.494
R231 vdd.n212 vdd.n190 190.494
R232 vdd.n203 vdd.n189 190.494
R233 vdd.n288 vdd.n254 190.494
R234 vdd.n280 vdd.n266 190.494
R235 vdd.n164 vdd.n143 190.494
R236 vdd.n171 vdd.n170 190.494
R237 vdd.n161 vdd.n160 190.494
R238 vdd.n156 vdd.n131 190.494
R239 vdd.n32 vdd.n19 179.118
R240 vdd.n33 vdd.n14 179.118
R241 vdd.n38 vdd.n14 179.118
R242 vdd.n40 vdd.n39 179.118
R243 vdd.n39 vdd.n11 179.118
R244 vdd.n49 vdd.n11 179.118
R245 vdd.n49 vdd.n6 179.118
R246 vdd.n80 vdd.n6 179.118
R247 vdd.n80 vdd.n79 179.118
R248 vdd.n78 vdd.n53 179.118
R249 vdd.n73 vdd.n53 179.118
R250 vdd.n72 vdd.n58 179.118
R251 vdd.n28 vdd.n27 173.642
R252 vdd.n68 vdd.n67 173.642
R253 vdd.n83 vdd.n2 131.388
R254 vdd.n51 vdd.n2 131.388
R255 vdd.n45 vdd.n44 131.388
R256 vdd.n45 vdd.n9 131.388
R257 vdd.n347 vdd.n178 131.388
R258 vdd.n352 vdd.n178 131.388
R259 vdd.n332 vdd.n230 131.388
R260 vdd.n333 vdd.n332 131.388
R261 vdd.n301 vdd.n252 131.388
R262 vdd.n321 vdd.n252 131.388
R263 vdd.n306 vdd.n293 131.388
R264 vdd.n307 vdd.n306 131.388
R265 vdd.n241 vdd.n240 131.388
R266 vdd.n245 vdd.n240 131.388
R267 vdd.n342 vdd.n341 131.388
R268 vdd.n341 vdd.n246 131.388
R269 vdd.n79 vdd.n78 120.168
R270 vdd.n33 vdd.n32 117.9
R271 vdd.n73 vdd.n72 117.9
R272 vdd vdd.n16 92.5005
R273 vdd.n16 vdd.n14 92.5005
R274 vdd.n18 vdd.n15 92.5005
R275 vdd.n15 vdd.n14 92.5005
R276 vdd.n52 vdd 92.5005
R277 vdd.n80 vdd.n52 92.5005
R278 vdd vdd.n50 92.5005
R279 vdd.n50 vdd.n49 92.5005
R280 vdd.n13 vdd 92.5005
R281 vdd.n39 vdd.n13 92.5005
R282 vdd.n43 vdd.n12 92.5005
R283 vdd.n39 vdd.n12 92.5005
R284 vdd.n48 vdd.n1 92.5005
R285 vdd.n49 vdd.n48 92.5005
R286 vdd.n82 vdd.n81 92.5005
R287 vdd.n81 vdd.n80 92.5005
R288 vdd vdd.n55 92.5005
R289 vdd.n55 vdd.n53 92.5005
R290 vdd.n56 vdd.n54 92.5005
R291 vdd.n54 vdd.n53 92.5005
R292 vdd vdd.n60 92.5005
R293 vdd.n61 vdd.n59 92.5005
R294 vdd.n59 vdd.n58 92.5005
R295 vdd vdd.n21 92.5005
R296 vdd.n21 vdd.n19 92.5005
R297 vdd.n26 vdd.n20 92.5005
R298 vdd.n103 vdd 92.5005
R299 vdd.n108 vdd.n103 92.5005
R300 vdd.n102 vdd.n101 92.5005
R301 vdd.n104 vdd.n102 92.5005
R302 vdd.n92 vdd.n90 92.5005
R303 vdd.n95 vdd.n92 92.5005
R304 vdd.n91 vdd 92.5005
R305 vdd.n93 vdd.n91 92.5005
R306 vdd.n122 vdd.n99 92.5005
R307 vdd.n99 vdd.n95 92.5005
R308 vdd vdd.n98 92.5005
R309 vdd.n98 vdd.n93 92.5005
R310 vdd vdd.n110 92.5005
R311 vdd.n110 vdd.n108 92.5005
R312 vdd.n111 vdd.n109 92.5005
R313 vdd.n109 vdd.n104 92.5005
R314 vdd vdd.n260 92.5005
R315 vdd.n260 vdd.n258 92.5005
R316 vdd.n261 vdd.n259 92.5005
R317 vdd.n259 vdd.n258 92.5005
R318 vdd vdd.n183 92.5005
R319 vdd.n349 vdd.n183 92.5005
R320 vdd vdd.n234 92.5005
R321 vdd.n345 vdd.n234 92.5005
R322 vdd.n338 vdd 92.5005
R323 vdd.n338 vdd.n337 92.5005
R324 vdd.n328 vdd.n237 92.5005
R325 vdd.n337 vdd.n328 92.5005
R326 vdd.n344 vdd.n343 92.5005
R327 vdd.n345 vdd.n344 92.5005
R328 vdd.n242 vdd.n227 92.5005
R329 vdd.n349 vdd.n227 92.5005
R330 vdd vdd.n200 92.5005
R331 vdd.n200 vdd.n185 92.5005
R332 vdd.n201 vdd.n199 92.5005
R333 vdd.n199 vdd.n185 92.5005
R334 vdd vdd.n197 92.5005
R335 vdd.n197 vdd.n195 92.5005
R336 vdd.n198 vdd.n196 92.5005
R337 vdd.n196 vdd.n195 92.5005
R338 vdd.n274 vdd.n269 92.5005
R339 vdd.n269 vdd.n262 92.5005
R340 vdd vdd.n268 92.5005
R341 vdd.n268 vdd.n262 92.5005
R342 vdd.n257 vdd.n255 92.5005
R343 vdd.n258 vdd.n257 92.5005
R344 vdd.n256 vdd 92.5005
R345 vdd.n258 vdd.n256 92.5005
R346 vdd.n322 vdd.n251 92.5005
R347 vdd.n251 vdd.n249 92.5005
R348 vdd.n296 vdd.n253 92.5005
R349 vdd.n303 vdd.n296 92.5005
R350 vdd.n308 vdd.n292 92.5005
R351 vdd.n292 vdd.n290 92.5005
R352 vdd vdd.n291 92.5005
R353 vdd.n291 vdd.n290 92.5005
R354 vdd.n302 vdd 92.5005
R355 vdd.n303 vdd.n302 92.5005
R356 vdd vdd.n250 92.5005
R357 vdd.n250 vdd.n249 92.5005
R358 vdd.n351 vdd.n350 92.5005
R359 vdd.n350 vdd.n349 92.5005
R360 vdd.n233 vdd.n177 92.5005
R361 vdd.n345 vdd.n233 92.5005
R362 vdd.n334 vdd.n327 92.5005
R363 vdd.n337 vdd.n327 92.5005
R364 vdd.n336 vdd 92.5005
R365 vdd.n337 vdd.n336 92.5005
R366 vdd vdd.n346 92.5005
R367 vdd.n346 vdd.n345 92.5005
R368 vdd.n348 vdd 92.5005
R369 vdd.n349 vdd.n348 92.5005
R370 vdd.n222 vdd.n187 92.5005
R371 vdd.n187 vdd.n185 92.5005
R372 vdd vdd.n186 92.5005
R373 vdd.n186 vdd.n185 92.5005
R374 vdd.n194 vdd.n192 92.5005
R375 vdd.n195 vdd.n194 92.5005
R376 vdd.n193 vdd 92.5005
R377 vdd.n195 vdd.n193 92.5005
R378 vdd vdd.n265 92.5005
R379 vdd.n265 vdd.n262 92.5005
R380 vdd.n267 vdd.n264 92.5005
R381 vdd.n264 vdd.n262 92.5005
R382 vdd.n146 vdd 92.5005
R383 vdd.n151 vdd.n146 92.5005
R384 vdd.n145 vdd.n144 92.5005
R385 vdd.n147 vdd.n145 92.5005
R386 vdd.n135 vdd.n133 92.5005
R387 vdd.n138 vdd.n135 92.5005
R388 vdd.n134 vdd 92.5005
R389 vdd.n136 vdd.n134 92.5005
R390 vdd.n165 vdd.n142 92.5005
R391 vdd.n142 vdd.n138 92.5005
R392 vdd vdd.n141 92.5005
R393 vdd.n141 vdd.n136 92.5005
R394 vdd vdd.n153 92.5005
R395 vdd.n153 vdd.n151 92.5005
R396 vdd.n154 vdd.n152 92.5005
R397 vdd.n152 vdd.n147 92.5005
R398 vdd.n125 vdd.n93 91.6935
R399 vdd.n125 vdd.n95 91.6935
R400 vdd.n115 vdd.n104 91.6935
R401 vdd.n115 vdd.n108 91.6935
R402 vdd.n168 vdd.n136 91.6935
R403 vdd.n168 vdd.n138 91.6935
R404 vdd.n158 vdd.n147 91.6935
R405 vdd.n158 vdd.n151 91.6935
R406 vdd.n277 vdd.n262 89.559
R407 vdd.n282 vdd.n262 89.559
R408 vdd.n285 vdd.n258 89.559
R409 vdd.n312 vdd.n258 89.559
R410 vdd.n311 vdd.n290 89.559
R411 vdd.n304 vdd.n290 89.559
R412 vdd.n304 vdd.n303 89.559
R413 vdd.n303 vdd.n297 89.559
R414 vdd.n297 vdd.n249 89.559
R415 vdd.n325 vdd.n249 89.559
R416 vdd.n337 vdd.n326 89.559
R417 vdd.n337 vdd.n232 89.559
R418 vdd.n345 vdd.n232 89.559
R419 vdd.n345 vdd.n182 89.559
R420 vdd.n349 vdd.n182 89.559
R421 vdd.n349 vdd.n226 89.559
R422 vdd.n225 vdd.n185 89.559
R423 vdd.n206 vdd.n185 89.559
R424 vdd.n209 vdd.n195 89.559
R425 vdd.n214 vdd.n195 89.559
R426 vdd.n67 vdd.n60 79.4196
R427 vdd.n27 vdd.n20 79.4196
R428 vdd.n312 vdd.n311 60.084
R429 vdd.n326 vdd.n325 60.084
R430 vdd.n226 vdd.n225 60.084
R431 vdd.n44 vdd.n43 59.4829
R432 vdd.n44 vdd.n1 59.4829
R433 vdd.n83 vdd.n82 59.4829
R434 vdd vdd.n9 59.4829
R435 vdd vdd.n9 59.4829
R436 vdd.n51 vdd 59.4829
R437 vdd vdd.n51 59.4829
R438 vdd vdd.n230 59.4829
R439 vdd vdd.n230 59.4829
R440 vdd.n347 vdd 59.4829
R441 vdd vdd.n347 59.4829
R442 vdd.n334 vdd.n333 59.4829
R443 vdd.n333 vdd.n177 59.4829
R444 vdd.n352 vdd.n351 59.4829
R445 vdd.n293 vdd 59.4829
R446 vdd vdd.n293 59.4829
R447 vdd vdd.n301 59.4829
R448 vdd.n301 vdd 59.4829
R449 vdd.n308 vdd.n307 59.4829
R450 vdd.n307 vdd.n253 59.4829
R451 vdd.n322 vdd.n321 59.4829
R452 vdd.n342 vdd.n237 59.4829
R453 vdd.n343 vdd.n342 59.4829
R454 vdd.n242 vdd.n241 59.4829
R455 vdd vdd.n246 59.4829
R456 vdd.n246 vdd 59.4829
R457 vdd vdd.n245 59.4829
R458 vdd.n245 vdd 59.4829
R459 vdd.n84 vdd.n83 59.1064
R460 vdd.n353 vdd.n352 59.1064
R461 vdd.n321 vdd.n320 59.1064
R462 vdd.n241 vdd.n175 59.1064
R463 vdd.n285 vdd.n282 58.9504
R464 vdd.n209 vdd.n206 58.9504
R465 vdd.n104 vdd.n95 26.5564
R466 vdd.n147 vdd.n138 26.5564
R467 vdd.n37 vdd.n36 23.1255
R468 vdd.n38 vdd.n37 23.1255
R469 vdd.n35 vdd.n34 23.1255
R470 vdd.n34 vdd.n33 23.1255
R471 vdd.n46 vdd.n45 23.1255
R472 vdd.n46 vdd.n11 23.1255
R473 vdd.n7 vdd.n2 23.1255
R474 vdd.n7 vdd.n6 23.1255
R475 vdd.n5 vdd.n3 23.1255
R476 vdd.n79 vdd.n5 23.1255
R477 vdd.n42 vdd.n41 23.1255
R478 vdd.n41 vdd.n40 23.1255
R479 vdd.n75 vdd.n74 23.1255
R480 vdd.n74 vdd.n73 23.1255
R481 vdd.n77 vdd.n76 23.1255
R482 vdd.n78 vdd.n77 23.1255
R483 vdd.n69 vdd.n68 23.1255
R484 vdd.n71 vdd.n70 23.1255
R485 vdd.n72 vdd.n71 23.1255
R486 vdd.n31 vdd.n30 23.1255
R487 vdd.n32 vdd.n31 23.1255
R488 vdd.n29 vdd.n28 23.1255
R489 vdd.n117 vdd.n116 23.1255
R490 vdd.n116 vdd.n115 23.1255
R491 vdd.n107 vdd.n106 23.1255
R492 vdd.n115 vdd.n107 23.1255
R493 vdd.n127 vdd.n126 23.1255
R494 vdd.n126 vdd.n125 23.1255
R495 vdd.n97 vdd.n96 23.1255
R496 vdd.n125 vdd.n97 23.1255
R497 vdd.n100 vdd.n94 23.1255
R498 vdd.n125 vdd.n94 23.1255
R499 vdd.n124 vdd.n123 23.1255
R500 vdd.n125 vdd.n124 23.1255
R501 vdd.n114 vdd.n113 23.1255
R502 vdd.n115 vdd.n114 23.1255
R503 vdd.n112 vdd.n105 23.1255
R504 vdd.n115 vdd.n105 23.1255
R505 vdd.n289 vdd.n288 23.1255
R506 vdd.n312 vdd.n289 23.1255
R507 vdd.n287 vdd.n286 23.1255
R508 vdd.n286 vdd.n285 23.1255
R509 vdd.n341 vdd.n340 23.1255
R510 vdd.n340 vdd.n232 23.1255
R511 vdd.n240 vdd.n239 23.1255
R512 vdd.n239 vdd.n182 23.1255
R513 vdd.n244 vdd.n243 23.1255
R514 vdd.n243 vdd.n226 23.1255
R515 vdd.n248 vdd.n247 23.1255
R516 vdd.n326 vdd.n247 23.1255
R517 vdd.n204 vdd.n203 23.1255
R518 vdd.n206 vdd.n204 23.1255
R519 vdd.n202 vdd.n184 23.1255
R520 vdd.n225 vdd.n184 23.1255
R521 vdd.n213 vdd.n212 23.1255
R522 vdd.n214 vdd.n213 23.1255
R523 vdd.n211 vdd.n210 23.1255
R524 vdd.n210 vdd.n209 23.1255
R525 vdd.n270 vdd.n263 23.1255
R526 vdd.n282 vdd.n263 23.1255
R527 vdd.n276 vdd.n275 23.1255
R528 vdd.n277 vdd.n276 23.1255
R529 vdd.n314 vdd.n313 23.1255
R530 vdd.n313 vdd.n312 23.1255
R531 vdd.n284 vdd.n283 23.1255
R532 vdd.n285 vdd.n284 23.1255
R533 vdd.n306 vdd.n305 23.1255
R534 vdd.n305 vdd.n304 23.1255
R535 vdd.n299 vdd.n252 23.1255
R536 vdd.n299 vdd.n297 23.1255
R537 vdd.n324 vdd.n323 23.1255
R538 vdd.n325 vdd.n324 23.1255
R539 vdd.n310 vdd.n309 23.1255
R540 vdd.n311 vdd.n310 23.1255
R541 vdd.n332 vdd.n331 23.1255
R542 vdd.n331 vdd.n232 23.1255
R543 vdd.n228 vdd.n178 23.1255
R544 vdd.n228 vdd.n182 23.1255
R545 vdd.n181 vdd.n179 23.1255
R546 vdd.n226 vdd.n181 23.1255
R547 vdd.n335 vdd.n329 23.1255
R548 vdd.n329 vdd.n326 23.1255
R549 vdd.n205 vdd.n188 23.1255
R550 vdd.n206 vdd.n205 23.1255
R551 vdd.n224 vdd.n223 23.1255
R552 vdd.n225 vdd.n224 23.1255
R553 vdd.n216 vdd.n215 23.1255
R554 vdd.n215 vdd.n214 23.1255
R555 vdd.n208 vdd.n207 23.1255
R556 vdd.n209 vdd.n208 23.1255
R557 vdd.n281 vdd.n280 23.1255
R558 vdd.n282 vdd.n281 23.1255
R559 vdd.n279 vdd.n278 23.1255
R560 vdd.n278 vdd.n277 23.1255
R561 vdd.n160 vdd.n159 23.1255
R562 vdd.n159 vdd.n158 23.1255
R563 vdd.n150 vdd.n149 23.1255
R564 vdd.n158 vdd.n150 23.1255
R565 vdd.n170 vdd.n169 23.1255
R566 vdd.n169 vdd.n168 23.1255
R567 vdd.n140 vdd.n139 23.1255
R568 vdd.n168 vdd.n140 23.1255
R569 vdd.n143 vdd.n137 23.1255
R570 vdd.n168 vdd.n137 23.1255
R571 vdd.n167 vdd.n166 23.1255
R572 vdd.n168 vdd.n167 23.1255
R573 vdd.n157 vdd.n156 23.1255
R574 vdd.n158 vdd.n157 23.1255
R575 vdd.n155 vdd.n148 23.1255
R576 vdd.n158 vdd.n148 23.1255
R577 vdd.n67 vdd.n58 8.97701
R578 vdd.n27 vdd.n19 8.97701
R579 vdd vdd.n86 2.79913
R580 vdd.n64 vdd 2.3405
R581 vdd.n63 vdd 2.3405
R582 vdd.n22 vdd 2.3405
R583 vdd.n24 vdd 2.3405
R584 vdd.n89 vdd 2.3405
R585 vdd.n89 vdd 2.3405
R586 vdd.n119 vdd 2.3405
R587 vdd.n119 vdd 2.3405
R588 vdd.n271 vdd 2.3405
R589 vdd.n271 vdd 2.3405
R590 vdd.n317 vdd 2.3405
R591 vdd.n317 vdd 2.3405
R592 vdd.n219 vdd 2.3405
R593 vdd.n219 vdd 2.3405
R594 vdd.n191 vdd 2.3405
R595 vdd.n191 vdd 2.3405
R596 vdd.n132 vdd 2.3405
R597 vdd.n132 vdd 2.3405
R598 vdd.n162 vdd 2.3405
R599 vdd.n162 vdd 2.3405
R600 vdd.n0 vdd 2.29412
R601 vdd.n318 vdd 2.29412
R602 vdd.n176 vdd 2.29412
R603 vdd.n176 vdd 2.29412
R604 vdd.n25 vdd.n24 2.07925
R605 vdd.n130 vdd.n87 2.02473
R606 vdd.n23 vdd.n17 1.8605
R607 vdd.n62 vdd.n57 1.8605
R608 vdd.n66 vdd.n65 1.8605
R609 vdd.n129 vdd.n88 1.8605
R610 vdd.n120 vdd.n118 1.8605
R611 vdd.n129 vdd.n128 1.8605
R612 vdd.n121 vdd.n120 1.8605
R613 vdd.n272 vdd.n266 1.8605
R614 vdd.n316 vdd.n254 1.8605
R615 vdd.n220 vdd.n189 1.8605
R616 vdd.n218 vdd.n190 1.8605
R617 vdd.n273 vdd.n272 1.8605
R618 vdd.n316 vdd.n315 1.8605
R619 vdd.n221 vdd.n220 1.8605
R620 vdd.n218 vdd.n217 1.8605
R621 vdd.n172 vdd.n131 1.8605
R622 vdd.n163 vdd.n161 1.8605
R623 vdd.n172 vdd.n171 1.8605
R624 vdd.n164 vdd.n163 1.8605
R625 vdd.n357 vdd.n356 1.76063
R626 vdd.n173 vdd.n87 1.75125
R627 vdd.n86 vdd 1.65831
R628 vdd.n356 vdd.n174 1.28995
R629 vdd.n174 vdd.n130 1.28887
R630 vdd.n174 vdd.n173 1.06531
R631 vdd.n130 vdd.n129 1.06168
R632 vdd.n173 vdd.n172 1.06168
R633 vdd.n86 vdd.n85 0.814562
R634 vdd.n85 vdd.n0 0.720812
R635 vdd.n85 vdd.n84 0.715885
R636 vdd.n354 vdd.n175 0.715885
R637 vdd.n320 vdd.n319 0.715885
R638 vdd.n354 vdd.n353 0.715885
R639 vdd.n319 vdd 0.413
R640 vdd.n355 vdd.n354 0.410656
R641 vdd.n66 vdd.n61 0.376971
R642 vdd.n57 vdd.n56 0.376971
R643 vdd.n84 vdd.n1 0.376971
R644 vdd.n18 vdd.n17 0.376971
R645 vdd.n26 vdd.n25 0.376971
R646 vdd.n122 vdd.n121 0.376971
R647 vdd.n128 vdd.n90 0.376971
R648 vdd.n118 vdd.n101 0.376971
R649 vdd.n111 vdd.n88 0.376971
R650 vdd.n217 vdd.n192 0.376971
R651 vdd.n222 vdd.n221 0.376971
R652 vdd.n353 vdd.n177 0.376971
R653 vdd.n320 vdd.n253 0.376971
R654 vdd.n315 vdd.n255 0.376971
R655 vdd.n274 vdd.n273 0.376971
R656 vdd.n198 vdd.n190 0.376971
R657 vdd.n201 vdd.n189 0.376971
R658 vdd.n343 vdd.n175 0.376971
R659 vdd.n261 vdd.n254 0.376971
R660 vdd.n267 vdd.n266 0.376971
R661 vdd.n165 vdd.n164 0.376971
R662 vdd.n171 vdd.n133 0.376971
R663 vdd.n161 vdd.n144 0.376971
R664 vdd.n154 vdd.n131 0.376971
R665 vdd.n319 vdd.n318 0.360656
R666 vdd.n354 vdd.n176 0.360656
R667 vdd.n62 vdd 0.33175
R668 vdd vdd.n23 0.328625
R669 vdd.n65 vdd 0.328625
R670 vdd.n357 vdd.n87 0.263158
R671 vdd.n23 vdd.n22 0.21925
R672 vdd.n63 vdd.n62 0.21925
R673 vdd.n65 vdd.n64 0.21925
R674 vdd.n220 vdd 0.166125
R675 vdd.n120 vdd 0.164562
R676 vdd.n316 vdd 0.164562
R677 vdd vdd.n218 0.164562
R678 vdd.n163 vdd 0.164562
R679 vdd.n24 vdd 0.109875
R680 vdd.n22 vdd 0.109875
R681 vdd vdd.n63 0.109875
R682 vdd.n64 vdd 0.109875
R683 vdd.n129 vdd.n89 0.109875
R684 vdd.n120 vdd.n119 0.109875
R685 vdd.n272 vdd.n271 0.109875
R686 vdd.n317 vdd.n316 0.109875
R687 vdd.n220 vdd.n219 0.109875
R688 vdd.n218 vdd.n191 0.109875
R689 vdd.n172 vdd.n132 0.109875
R690 vdd.n163 vdd.n162 0.109875
R691 vdd vdd.n0 0.102062
R692 vdd.n356 vdd.n355 0.0780862
R693 vdd vdd.n89 0.0551875
R694 vdd.n119 vdd 0.0551875
R695 vdd.n271 vdd 0.0551875
R696 vdd vdd.n317 0.0551875
R697 vdd.n219 vdd 0.0551875
R698 vdd.n191 vdd 0.0551875
R699 vdd vdd.n132 0.0551875
R700 vdd.n162 vdd 0.0551875
R701 vdd.n318 vdd 0.0512812
R702 vdd vdd.n176 0.0512812
R703 vdd vdd.n357 0.00538077
R704 vdd.n355 vdd 0.00284375
R705 vss.n107 vss.n106 4116.13
R706 vss.n298 vss.n207 2547.63
R707 vss.n203 vss.n187 2510.19
R708 vss.n306 vss.n202 2306.06
R709 vss.n306 vss.n203 2306.06
R710 vss.n202 vss.n187 2306.06
R711 vss.n234 vss.n201 2306.06
R712 vss.n237 vss.n201 2306.06
R713 vss.n234 vss.n185 2306.06
R714 vss.n237 vss.n185 2306.06
R715 vss.n323 vss.n308 2306.06
R716 vss.n308 vss.n189 2306.06
R717 vss.n314 vss.n307 2306.06
R718 vss.n314 vss.n188 2306.06
R719 vss.n327 vss.n199 2306.06
R720 vss.n328 vss.n327 2306.06
R721 vss.n199 vss.n184 2306.06
R722 vss.n328 vss.n184 2306.06
R723 vss.n325 vss.n190 2306.06
R724 vss.n325 vss.n191 2306.06
R725 vss.n335 vss.n190 2306.06
R726 vss.n335 vss.n191 2306.06
R727 vss.n220 vss.n207 2306.06
R728 vss.n220 vss.n208 2306.06
R729 vss.n298 vss.n208 2306.06
R730 vss.n232 vss.n218 2306.06
R731 vss.n245 vss.n232 2306.06
R732 vss.n233 vss.n218 2306.06
R733 vss.n245 vss.n233 2306.06
R734 vss.n247 vss.n216 2306.06
R735 vss.n252 vss.n216 2306.06
R736 vss.n260 vss.n246 2306.06
R737 vss.n264 vss.n246 2306.06
R738 vss.n221 vss.n212 2306.06
R739 vss.n221 vss.n213 2306.06
R740 vss.n225 vss.n212 2306.06
R741 vss.n225 vss.n213 2306.06
R742 vss.n226 vss.n210 2306.06
R743 vss.n226 vss.n211 2306.06
R744 vss.n230 vss.n210 2306.06
R745 vss.n230 vss.n211 2306.06
R746 vss.n275 vss.n214 2306.06
R747 vss.n277 vss.n214 2306.06
R748 vss.n287 vss.n271 2306.06
R749 vss.n290 vss.n271 2306.06
R750 vss.n153 vss.n135 2306.06
R751 vss.n144 vss.n135 2306.06
R752 vss.n153 vss.n136 2306.06
R753 vss.n144 vss.n136 2306.06
R754 vss.n125 vss.n120 2306.06
R755 vss.n132 vss.n125 2306.06
R756 vss.n126 vss.n120 2306.06
R757 vss.n132 vss.n126 2306.06
R758 vss.n110 vss.n81 2306.06
R759 vss.n108 vss.n81 2306.06
R760 vss.n164 vss.n118 2306.06
R761 vss.n119 vss.n118 2306.06
R762 vss.n94 vss.n83 2306.06
R763 vss.n105 vss.n83 2306.06
R764 vss.n94 vss.n84 2306.06
R765 vss.n105 vss.n84 2306.06
R766 vss.n97 vss.n87 2306.06
R767 vss.n90 vss.n88 2306.06
R768 vss.n97 vss.n88 2306.06
R769 vss.n142 vss.n133 2306.06
R770 vss.n146 vss.n142 2306.06
R771 vss.n143 vss.n133 2306.06
R772 vss.n146 vss.n143 2306.06
R773 vss.n160 vss.n122 2306.06
R774 vss.n156 vss.n122 2306.06
R775 vss.n160 vss.n123 2306.06
R776 vss.n156 vss.n123 2306.06
R777 vss.n62 vss.n36 2306.06
R778 vss.n36 vss.n32 2306.06
R779 vss.n62 vss.n37 2306.06
R780 vss.n37 vss.n32 2306.06
R781 vss.n35 vss.n29 2306.06
R782 vss.n64 vss.n29 2306.06
R783 vss.n35 vss.n30 2306.06
R784 vss.n64 vss.n30 2306.06
R785 vss.n46 vss.n41 2306.06
R786 vss.n55 vss.n41 2306.06
R787 vss.n46 vss.n42 2306.06
R788 vss.n55 vss.n42 2306.06
R789 vss.n48 vss.n44 2306.06
R790 vss.n53 vss.n48 2306.06
R791 vss.n49 vss.n44 2306.06
R792 vss.n53 vss.n49 2306.06
R793 vss.n19 vss.n9 2306.06
R794 vss.n13 vss.n9 2306.06
R795 vss.n19 vss.n10 2306.06
R796 vss.n22 vss.n2 2306.06
R797 vss.n22 vss.n3 2306.06
R798 vss.n5 vss.n3 2306.06
R799 vss.n312 vss.n311 1390.59
R800 vss.n312 vss.n182 1390.59
R801 vss.n319 vss.n309 1390.59
R802 vss.n319 vss.n181 1390.59
R803 vss.n259 vss.n217 1390.59
R804 vss.n265 vss.n217 1390.59
R805 vss.n270 vss.n248 1390.59
R806 vss.n270 vss.n249 1390.59
R807 vss.n296 vss.n272 1390.59
R808 vss.n296 vss.n273 1390.59
R809 vss.n286 vss.n215 1390.59
R810 vss.n291 vss.n215 1390.59
R811 vss.n115 vss.n79 1390.59
R812 vss.n115 vss.n75 1390.59
R813 vss.n112 vss.n78 1390.59
R814 vss.n112 vss.n74 1390.59
R815 vss.n21 vss.n7 1121.29
R816 vss.n20 vss.n8 1121.29
R817 vss.n323 vss.n309 915.471
R818 vss.n309 vss.n200 915.471
R819 vss.n311 vss.n200 915.471
R820 vss.n311 vss.n307 915.471
R821 vss.n189 vss.n181 915.471
R822 vss.n337 vss.n181 915.471
R823 vss.n337 vss.n182 915.471
R824 vss.n188 vss.n182 915.471
R825 vss.n248 vss.n247 915.471
R826 vss.n258 vss.n248 915.471
R827 vss.n259 vss.n258 915.471
R828 vss.n260 vss.n259 915.471
R829 vss.n252 vss.n249 915.471
R830 vss.n266 vss.n249 915.471
R831 vss.n266 vss.n265 915.471
R832 vss.n265 vss.n264 915.471
R833 vss.n275 vss.n272 915.471
R834 vss.n285 vss.n272 915.471
R835 vss.n286 vss.n285 915.471
R836 vss.n287 vss.n286 915.471
R837 vss.n277 vss.n273 915.471
R838 vss.n292 vss.n273 915.471
R839 vss.n292 vss.n291 915.471
R840 vss.n291 vss.n290 915.471
R841 vss.n110 vss.n78 915.471
R842 vss.n168 vss.n78 915.471
R843 vss.n168 vss.n79 915.471
R844 vss.n164 vss.n79 915.471
R845 vss.n108 vss.n74 915.471
R846 vss.n170 vss.n74 915.471
R847 vss.n170 vss.n75 915.471
R848 vss.n119 vss.n75 915.471
R849 vss.n6 vss.n5 744.25
R850 vss.n13 vss.n12 744.25
R851 vss.n21 vss.n20 738.066
R852 vss.n96 vss.n92 560.645
R853 vss.n95 vss.n82 560.645
R854 vss.n106 vss.n82 560.645
R855 vss.n109 vss.n107 560.645
R856 vss.n109 vss.n76 560.645
R857 vss.n169 vss.n76 560.645
R858 vss.n169 vss.n77 560.645
R859 vss.n163 vss.n77 560.645
R860 vss.n163 vss.n162 560.645
R861 vss.n161 vss.n121 560.645
R862 vss.n155 vss.n121 560.645
R863 vss.n154 vss.n134 560.645
R864 vss.n145 vss.n134 560.645
R865 vss.n91 vss.n90 476.983
R866 vss.n162 vss.n161 376.13
R867 vss.n96 vss.n95 369.033
R868 vss.n155 vss.n154 369.033
R869 vss.n251 vss.n250 343.154
R870 vss.n326 vss.n183 298.207
R871 vss.n336 vss.n183 298.207
R872 vss.n297 vss.n209 298.207
R873 vss.n297 vss.n231 298.207
R874 vss.n63 vss.n31 298.207
R875 vss.n63 vss.n33 298.207
R876 vss.n54 vss.n43 298.207
R877 vss.n54 vss.n47 298.207
R878 vss.n230 vss.n229 292.5
R879 vss.n231 vss.n230 292.5
R880 vss vss.n226 292.5
R881 vss.n226 vss.n209 292.5
R882 vss.n225 vss.n224 292.5
R883 vss.n231 vss.n225 292.5
R884 vss vss.n221 292.5
R885 vss.n221 vss.n209 292.5
R886 vss.n264 vss.n263 292.5
R887 vss.n264 vss.n231 292.5
R888 vss.n267 vss.n266 292.5
R889 vss.n266 vss.n231 292.5
R890 vss.n253 vss.n252 292.5
R891 vss.n252 vss.n231 292.5
R892 vss.n247 vss 292.5
R893 vss.n247 vss.n209 292.5
R894 vss.n258 vss 292.5
R895 vss.n258 vss.n209 292.5
R896 vss vss.n260 292.5
R897 vss.n260 vss.n209 292.5
R898 vss.n243 vss.n233 292.5
R899 vss.n233 vss.n231 292.5
R900 vss vss.n232 292.5
R901 vss.n232 vss.n209 292.5
R902 vss.n208 vss.n206 292.5
R903 vss.n231 vss.n208 292.5
R904 vss.n207 vss 292.5
R905 vss.n209 vss.n207 292.5
R906 vss.n335 vss 292.5
R907 vss.n336 vss.n335 292.5
R908 vss.n325 vss.n324 292.5
R909 vss.n326 vss.n325 292.5
R910 vss vss.n184 292.5
R911 vss.n336 vss.n184 292.5
R912 vss.n327 vss.n197 292.5
R913 vss.n327 vss.n326 292.5
R914 vss vss.n188 292.5
R915 vss.n336 vss.n188 292.5
R916 vss vss.n337 292.5
R917 vss.n337 vss.n336 292.5
R918 vss vss.n189 292.5
R919 vss.n336 vss.n189 292.5
R920 vss.n323 vss.n322 292.5
R921 vss.n326 vss.n323 292.5
R922 vss.n318 vss.n200 292.5
R923 vss.n326 vss.n200 292.5
R924 vss.n316 vss.n307 292.5
R925 vss.n326 vss.n307 292.5
R926 vss vss.n185 292.5
R927 vss.n336 vss.n185 292.5
R928 vss.n236 vss.n201 292.5
R929 vss.n326 vss.n201 292.5
R930 vss vss.n187 292.5
R931 vss.n336 vss.n187 292.5
R932 vss.n306 vss.n305 292.5
R933 vss.n326 vss.n306 292.5
R934 vss.n290 vss.n289 292.5
R935 vss.n290 vss.n231 292.5
R936 vss.n293 vss.n292 292.5
R937 vss.n292 vss.n231 292.5
R938 vss.n278 vss.n277 292.5
R939 vss.n277 vss.n231 292.5
R940 vss vss.n275 292.5
R941 vss.n275 vss.n209 292.5
R942 vss.n285 vss 292.5
R943 vss.n285 vss.n209 292.5
R944 vss vss.n287 292.5
R945 vss.n287 vss.n209 292.5
R946 vss.n143 vss.n141 292.5
R947 vss.n143 vss.n134 292.5
R948 vss.n142 vss 292.5
R949 vss.n142 vss.n134 292.5
R950 vss.n88 vss 292.5
R951 vss.n92 vss.n88 292.5
R952 vss.n87 vss.n86 292.5
R953 vss vss.n84 292.5
R954 vss.n84 vss.n82 292.5
R955 vss.n85 vss.n83 292.5
R956 vss.n83 vss.n82 292.5
R957 vss.n119 vss 292.5
R958 vss.n163 vss.n119 292.5
R959 vss vss.n170 292.5
R960 vss.n170 vss.n169 292.5
R961 vss.n108 vss 292.5
R962 vss.n109 vss.n108 292.5
R963 vss.n111 vss.n110 292.5
R964 vss.n110 vss.n109 292.5
R965 vss.n168 vss.n167 292.5
R966 vss.n169 vss.n168 292.5
R967 vss.n165 vss.n164 292.5
R968 vss.n164 vss.n163 292.5
R969 vss vss.n126 292.5
R970 vss.n126 vss.n121 292.5
R971 vss.n127 vss.n125 292.5
R972 vss.n125 vss.n121 292.5
R973 vss vss.n136 292.5
R974 vss.n136 vss.n134 292.5
R975 vss.n137 vss.n135 292.5
R976 vss.n135 vss.n134 292.5
R977 vss.n158 vss.n123 292.5
R978 vss.n123 vss.n121 292.5
R979 vss vss.n122 292.5
R980 vss.n122 vss.n121 292.5
R981 vss.n42 vss.n40 292.5
R982 vss.n47 vss.n42 292.5
R983 vss.n41 vss 292.5
R984 vss.n43 vss.n41 292.5
R985 vss.n30 vss 292.5
R986 vss.n33 vss.n30 292.5
R987 vss.n29 vss.n28 292.5
R988 vss.n31 vss.n29 292.5
R989 vss vss.n37 292.5
R990 vss.n37 vss.n33 292.5
R991 vss.n38 vss.n36 292.5
R992 vss.n36 vss.n31 292.5
R993 vss.n51 vss.n49 292.5
R994 vss.n49 vss.n47 292.5
R995 vss vss.n48 292.5
R996 vss.n48 vss.n43 292.5
R997 vss vss.n10 292.5
R998 vss.n11 vss.n9 292.5
R999 vss.n9 vss.n8 292.5
R1000 vss.n2 vss.n1 292.5
R1001 vss.n3 vss 292.5
R1002 vss.n7 vss.n3 292.5
R1003 vss.n261 vss.n256 249.667
R1004 vss.n91 vss.n87 205.887
R1005 vss.n12 vss.n10 175.803
R1006 vss.n6 vss.n2 175.803
R1007 vss.n289 vss.n288 150.418
R1008 vss.n316 vss.n315 150.417
R1009 vss.n263 vss.n262 150.417
R1010 vss.n165 vss.n117 150.417
R1011 vss.n305 vss.n204 149.835
R1012 vss.n305 vss.n304 149.835
R1013 vss vss.n204 149.835
R1014 vss.n236 vss.n235 149.835
R1015 vss.n238 vss.n236 149.835
R1016 vss.n235 vss 149.835
R1017 vss.n322 vss.n310 149.835
R1018 vss.n198 vss.n197 149.835
R1019 vss.n329 vss.n197 149.835
R1020 vss.n198 vss 149.835
R1021 vss.n324 vss.n192 149.835
R1022 vss.n324 vss.n193 149.835
R1023 vss vss.n192 149.835
R1024 vss.n219 vss 149.835
R1025 vss.n219 vss.n206 149.835
R1026 vss.n299 vss.n206 149.835
R1027 vss.n242 vss 149.835
R1028 vss.n243 vss.n242 149.835
R1029 vss.n244 vss.n243 149.835
R1030 vss.n253 vss.n251 149.835
R1031 vss.n222 vss 149.835
R1032 vss.n224 vss.n222 149.835
R1033 vss.n224 vss.n223 149.835
R1034 vss.n227 vss 149.835
R1035 vss.n229 vss.n227 149.835
R1036 vss.n229 vss.n228 149.835
R1037 vss.n278 vss.n276 149.835
R1038 vss.n152 vss.n137 149.835
R1039 vss.n138 vss.n137 149.835
R1040 vss.n152 vss 149.835
R1041 vss.n128 vss.n127 149.835
R1042 vss.n131 vss.n127 149.835
R1043 vss vss.n128 149.835
R1044 vss.n111 vss.n80 149.835
R1045 vss.n93 vss.n85 149.835
R1046 vss.n104 vss.n85 149.835
R1047 vss.n93 vss 149.835
R1048 vss.n89 vss.n86 149.835
R1049 vss.n98 vss.n86 149.835
R1050 vss.n89 vss 149.835
R1051 vss.n140 vss 149.835
R1052 vss.n141 vss.n140 149.835
R1053 vss.n147 vss.n141 149.835
R1054 vss.n158 vss.n157 149.835
R1055 vss.n159 vss.n158 149.835
R1056 vss.n159 vss 149.835
R1057 vss.n61 vss.n38 149.835
R1058 vss.n39 vss.n38 149.835
R1059 vss.n61 vss 149.835
R1060 vss.n34 vss.n28 149.835
R1061 vss.n65 vss.n28 149.835
R1062 vss.n34 vss 149.835
R1063 vss.n45 vss 149.835
R1064 vss.n45 vss.n40 149.835
R1065 vss.n56 vss.n40 149.835
R1066 vss.n52 vss.n51 149.835
R1067 vss.n51 vss.n50 149.835
R1068 vss.n50 vss 149.835
R1069 vss.n18 vss.n11 149.835
R1070 vss.n14 vss.n11 149.835
R1071 vss.n18 vss 149.835
R1072 vss.n4 vss.n1 149.835
R1073 vss.n4 vss 149.835
R1074 vss.n23 vss.n1 149.835
R1075 vss.n304 vss.n303 149.459
R1076 vss.n239 vss.n238 149.459
R1077 vss.n330 vss.n329 149.459
R1078 vss.n334 vss.n193 149.459
R1079 vss.n300 vss.n299 149.459
R1080 vss.n244 vss.n241 149.459
R1081 vss.n223 vss.n195 149.459
R1082 vss.n228 vss.n194 149.459
R1083 vss.n151 vss.n138 149.459
R1084 vss.n131 vss.n130 149.459
R1085 vss.n104 vss.n103 149.459
R1086 vss.n99 vss.n98 149.459
R1087 vss.n148 vss.n147 149.459
R1088 vss.n157 vss.n124 149.459
R1089 vss.n60 vss.n39 149.459
R1090 vss.n66 vss.n65 149.459
R1091 vss.n57 vss.n56 149.459
R1092 vss.n52 vss.n27 149.459
R1093 vss.n17 vss.n14 149.459
R1094 vss.n24 vss.n23 149.459
R1095 vss.n257 vss.n256 132.8
R1096 vss.n288 vss 132.129
R1097 vss.n315 vss 132.127
R1098 vss vss.n117 132.127
R1099 vss.n310 vss 130.802
R1100 vss.n276 vss 130.802
R1101 vss vss.n80 130.802
R1102 vss.n43 vss.n33 122.996
R1103 vss.n257 vss.n250 120.001
R1104 vss vss 118.966
R1105 vss.n228 vss.n211 117.001
R1106 vss.n297 vss.n211 117.001
R1107 vss.n227 vss.n210 117.001
R1108 vss.n297 vss.n210 117.001
R1109 vss.n223 vss.n213 117.001
R1110 vss.n297 vss.n213 117.001
R1111 vss.n222 vss.n212 117.001
R1112 vss.n297 vss.n212 117.001
R1113 vss.n270 vss.n269 117.001
R1114 vss.n297 vss.n270 117.001
R1115 vss.n255 vss.n217 117.001
R1116 vss.n297 vss.n217 117.001
R1117 vss.n262 vss.n246 117.001
R1118 vss.n297 vss.n246 117.001
R1119 vss.n251 vss.n216 117.001
R1120 vss.n297 vss.n216 117.001
R1121 vss.n245 vss.n244 117.001
R1122 vss.n297 vss.n245 117.001
R1123 vss.n242 vss.n218 117.001
R1124 vss.n297 vss.n218 117.001
R1125 vss.n299 vss.n298 117.001
R1126 vss.n298 vss.n297 117.001
R1127 vss.n220 vss.n219 117.001
R1128 vss.n297 vss.n220 117.001
R1129 vss.n193 vss.n191 117.001
R1130 vss.n191 vss.n183 117.001
R1131 vss.n192 vss.n190 117.001
R1132 vss.n190 vss.n183 117.001
R1133 vss.n329 vss.n328 117.001
R1134 vss.n328 vss.n183 117.001
R1135 vss.n199 vss.n198 117.001
R1136 vss.n199 vss.n183 117.001
R1137 vss.n320 vss.n319 117.001
R1138 vss.n319 vss.n183 117.001
R1139 vss.n313 vss.n312 117.001
R1140 vss.n312 vss.n183 117.001
R1141 vss.n315 vss.n314 117.001
R1142 vss.n314 vss.n183 117.001
R1143 vss.n310 vss.n308 117.001
R1144 vss.n308 vss.n183 117.001
R1145 vss.n238 vss.n237 117.001
R1146 vss.n237 vss.n183 117.001
R1147 vss.n235 vss.n234 117.001
R1148 vss.n234 vss.n183 117.001
R1149 vss.n304 vss.n203 117.001
R1150 vss.n203 vss.n183 117.001
R1151 vss.n204 vss.n202 117.001
R1152 vss.n202 vss.n183 117.001
R1153 vss.n296 vss.n295 117.001
R1154 vss.n297 vss.n296 117.001
R1155 vss.n280 vss.n215 117.001
R1156 vss.n297 vss.n215 117.001
R1157 vss.n288 vss.n271 117.001
R1158 vss.n297 vss.n271 117.001
R1159 vss.n276 vss.n214 117.001
R1160 vss.n297 vss.n214 117.001
R1161 vss.n147 vss.n146 117.001
R1162 vss.n146 vss.n145 117.001
R1163 vss.n140 vss.n133 117.001
R1164 vss.n154 vss.n133 117.001
R1165 vss.n98 vss.n97 117.001
R1166 vss.n97 vss.n96 117.001
R1167 vss.n90 vss.n89 117.001
R1168 vss.n105 vss.n104 117.001
R1169 vss.n106 vss.n105 117.001
R1170 vss.n94 vss.n93 117.001
R1171 vss.n95 vss.n94 117.001
R1172 vss.n113 vss.n112 117.001
R1173 vss.n112 vss.n76 117.001
R1174 vss.n116 vss.n115 117.001
R1175 vss.n115 vss.n77 117.001
R1176 vss.n118 vss.n117 117.001
R1177 vss.n162 vss.n118 117.001
R1178 vss.n81 vss.n80 117.001
R1179 vss.n107 vss.n81 117.001
R1180 vss.n132 vss.n131 117.001
R1181 vss.n155 vss.n132 117.001
R1182 vss.n128 vss.n120 117.001
R1183 vss.n161 vss.n120 117.001
R1184 vss.n144 vss.n138 117.001
R1185 vss.n145 vss.n144 117.001
R1186 vss.n153 vss.n152 117.001
R1187 vss.n154 vss.n153 117.001
R1188 vss.n157 vss.n156 117.001
R1189 vss.n156 vss.n155 117.001
R1190 vss.n160 vss.n159 117.001
R1191 vss.n161 vss.n160 117.001
R1192 vss.n56 vss.n55 117.001
R1193 vss.n55 vss.n54 117.001
R1194 vss.n46 vss.n45 117.001
R1195 vss.n54 vss.n46 117.001
R1196 vss.n65 vss.n64 117.001
R1197 vss.n64 vss.n63 117.001
R1198 vss.n35 vss.n34 117.001
R1199 vss.n63 vss.n35 117.001
R1200 vss.n39 vss.n32 117.001
R1201 vss.n63 vss.n32 117.001
R1202 vss.n62 vss.n61 117.001
R1203 vss.n63 vss.n62 117.001
R1204 vss.n53 vss.n52 117.001
R1205 vss.n54 vss.n53 117.001
R1206 vss.n50 vss.n44 117.001
R1207 vss.n54 vss.n44 117.001
R1208 vss.n14 vss.n13 117.001
R1209 vss.n19 vss.n18 117.001
R1210 vss.n20 vss.n19 117.001
R1211 vss.n5 vss.n4 117.001
R1212 vss.n23 vss.n22 117.001
R1213 vss.n22 vss.n21 117.001
R1214 vss vss.n177 115.576
R1215 vss.n12 vss.n8 94.4014
R1216 vss.n7 vss.n6 94.4014
R1217 vss.n281 vss.n280 90.3534
R1218 vss.n280 vss.n279 90.3534
R1219 vss.n317 vss.n313 90.3534
R1220 vss.n313 vss.n180 90.3534
R1221 vss.n321 vss.n320 90.3534
R1222 vss.n320 vss.n179 90.3534
R1223 vss.n256 vss.n255 90.3534
R1224 vss.n255 vss.n254 90.3534
R1225 vss.n269 vss.n250 90.3534
R1226 vss.n269 vss.n268 90.3534
R1227 vss.n295 vss.n274 90.3534
R1228 vss.n295 vss.n294 90.3534
R1229 vss.n166 vss.n116 90.3534
R1230 vss.n116 vss.n73 90.3534
R1231 vss.n114 vss.n113 90.3534
R1232 vss.n113 vss.n72 90.3534
R1233 vss.n262 vss.n261 89.9911
R1234 vss.n261 vss 77.2563
R1235 vss.n336 vss.n186 63.8191
R1236 vss.n92 vss.n91 60.5013
R1237 vss.n322 vss.n321 59.4829
R1238 vss.n321 vss.n318 59.4829
R1239 vss.n318 vss.n317 59.4829
R1240 vss.n317 vss.n316 59.4829
R1241 vss.n268 vss.n253 59.4829
R1242 vss.n268 vss.n267 59.4829
R1243 vss.n267 vss.n254 59.4829
R1244 vss.n263 vss.n254 59.4829
R1245 vss.n294 vss.n278 59.4829
R1246 vss.n294 vss.n293 59.4829
R1247 vss.n293 vss.n279 59.4829
R1248 vss.n289 vss.n279 59.4829
R1249 vss.n114 vss.n111 59.4829
R1250 vss.n167 vss.n114 59.4829
R1251 vss.n167 vss.n166 59.4829
R1252 vss.n166 vss.n165 59.4829
R1253 vss.n209 vss.n186 59.1777
R1254 vss vss.n179 40.4485
R1255 vss vss.n180 40.4485
R1256 vss vss.n180 40.4485
R1257 vss vss.n274 40.4485
R1258 vss vss.n281 40.4485
R1259 vss vss.n281 40.4485
R1260 vss vss.n72 40.4485
R1261 vss vss.n73 40.4485
R1262 vss vss.n73 40.4485
R1263 vss.n338 vss.n179 38.1445
R1264 vss.n284 vss.n274 38.1445
R1265 vss.n171 vss.n72 38.1445
R1266 vss.n174 vss.n70 5.57862
R1267 vss.n341 vss.n176 5.57706
R1268 vss.n178 vss 5.02361
R1269 vss.n178 vss 5.02361
R1270 vss.n282 vss 5.02361
R1271 vss.n71 vss 5.02361
R1272 vss.n332 vss 5.01717
R1273 vss.n332 vss 5.01717
R1274 vss.n196 vss 5.01717
R1275 vss.n196 vss 5.01717
R1276 vss.n205 vss 5.01717
R1277 vss.n205 vss 5.01717
R1278 vss.n301 vss 5.01717
R1279 vss.n301 vss 5.01717
R1280 vss.n100 vss 5.01717
R1281 vss.n101 vss 5.01717
R1282 vss.n139 vss 5.01717
R1283 vss.n139 vss 5.01717
R1284 vss.n149 vss 5.01717
R1285 vss.n149 vss 5.01717
R1286 vss.n26 vss 5.01717
R1287 vss.n26 vss 5.01717
R1288 vss.n58 vss 5.01717
R1289 vss.n58 vss 5.01717
R1290 vss.n0 vss 5.01717
R1291 vss.n15 vss 5.01717
R1292 vss.n69 vss.n25 4.58332
R1293 vss vss.n257 3.01226
R1294 vss.n69 vss.n68 2.46929
R1295 vss.n338 vss 2.3045
R1296 vss vss.n284 2.3045
R1297 vss.n171 vss 2.3045
R1298 vss.n100 vss.n99 1.96988
R1299 vss.n25 vss.n24 1.90103
R1300 vss.n333 vss.n194 1.8605
R1301 vss.n331 vss.n195 1.8605
R1302 vss.n241 vss.n240 1.8605
R1303 vss.n302 vss.n300 1.8605
R1304 vss.n334 vss.n333 1.8605
R1305 vss.n331 vss.n330 1.8605
R1306 vss.n240 vss.n239 1.8605
R1307 vss.n303 vss.n302 1.8605
R1308 vss.n129 vss.n124 1.8605
R1309 vss.n150 vss.n148 1.8605
R1310 vss.n103 vss.n102 1.8605
R1311 vss.n130 vss.n129 1.8605
R1312 vss.n151 vss.n150 1.8605
R1313 vss.n67 vss.n27 1.8605
R1314 vss.n59 vss.n57 1.8605
R1315 vss.n67 vss.n66 1.8605
R1316 vss.n60 vss.n59 1.8605
R1317 vss.n17 vss.n16 1.8605
R1318 vss.n342 vss.n341 1.79344
R1319 vss.n175 vss.n174 1.68993
R1320 vss.n173 vss 0.827844
R1321 vss.n284 vss.n283 0.715885
R1322 vss.n339 vss.n177 0.715885
R1323 vss.n339 vss.n338 0.715885
R1324 vss.n172 vss.n171 0.715885
R1325 vss.n283 vss 0.405187
R1326 vss.n340 vss.n339 0.402844
R1327 vss.n173 vss.n172 0.401281
R1328 vss.n303 vss 0.376971
R1329 vss.n239 vss 0.376971
R1330 vss.n330 vss 0.376971
R1331 vss vss.n334 0.376971
R1332 vss.n300 vss 0.376971
R1333 vss vss.n241 0.376971
R1334 vss.n257 vss.n177 0.376971
R1335 vss vss.n195 0.376971
R1336 vss vss.n194 0.376971
R1337 vss vss.n151 0.376971
R1338 vss.n130 vss 0.376971
R1339 vss.n103 vss 0.376971
R1340 vss.n99 vss 0.376971
R1341 vss.n148 vss 0.376971
R1342 vss.n124 vss 0.376971
R1343 vss vss.n60 0.376971
R1344 vss.n66 vss 0.376971
R1345 vss.n57 vss 0.376971
R1346 vss vss.n27 0.376971
R1347 vss vss.n17 0.376971
R1348 vss.n24 vss 0.376971
R1349 vss.n283 vss.n282 0.376281
R1350 vss.n339 vss.n178 0.376281
R1351 vss.n172 vss.n71 0.376281
R1352 vss.n16 vss 0.328625
R1353 vss.n342 vss.n175 0.250766
R1354 vss.n175 vss.n69 0.250595
R1355 vss.n16 vss.n15 0.21925
R1356 vss.n25 vss.n0 0.176322
R1357 vss.n240 vss 0.166125
R1358 vss.n129 vss 0.166125
R1359 vss vss.n331 0.164562
R1360 vss.n302 vss 0.164562
R1361 vss.n102 vss 0.164562
R1362 vss.n150 vss 0.164562
R1363 vss.n59 vss 0.164562
R1364 vss.n333 vss.n332 0.109875
R1365 vss.n331 vss.n196 0.109875
R1366 vss.n302 vss.n301 0.109875
R1367 vss.n102 vss.n101 0.109875
R1368 vss.n150 vss.n149 0.109875
R1369 vss.n59 vss.n58 0.109875
R1370 vss vss.n0 0.109875
R1371 vss.n15 vss 0.109875
R1372 vss.n129 vss.n70 0.0934687
R1373 vss.n240 vss.n176 0.0903438
R1374 vss.n68 vss.n26 0.0860255
R1375 vss.n341 vss.n340 0.0780862
R1376 vss.n174 vss.n173 0.0780862
R1377 vss.n332 vss 0.0551875
R1378 vss vss.n196 0.0551875
R1379 vss vss.n205 0.0551875
R1380 vss.n301 vss 0.0551875
R1381 vss vss.n100 0.0551875
R1382 vss.n101 vss 0.0551875
R1383 vss vss.n139 0.0551875
R1384 vss.n149 vss 0.0551875
R1385 vss vss.n26 0.0551875
R1386 vss.n58 vss 0.0551875
R1387 vss.n282 vss 0.0434688
R1388 vss vss.n178 0.0434688
R1389 vss vss.n71 0.0434688
R1390 vss.n68 vss.n67 0.0233551
R1391 vss.n205 vss.n176 0.0200312
R1392 vss.n139 vss.n70 0.0169062
R1393 vss vss.n342 0.00513139
R1394 vss.n340 vss 0.00284375
R1395 d0.n0 d0.t1 556.78
R1396 d0.t1 d0 547.24
R1397 d0 d0.t0 372.113
R1398 d0.n0 d0 9.54008
R1399 d0 d0.n0 0.141125
R1400 d0 d0 0.1255
R1401 d0 d0 0.063
R1402 d1.n0 d1.t1 556.78
R1403 d1.t1 d1 547.24
R1404 d1 d1.t0 372.113
R1405 d1.n0 d1 9.54008
R1406 d1 d1.n0 0.141125
R1407 d1 d1 0.1255
R1408 d1 d1 0.063
R1409 d2.n0 d2.t1 556.78
R1410 d2.t1 d2 547.24
R1411 d2 d2.t0 372.113
R1412 d2.n0 d2 9.54008
R1413 d2 d2.n0 0.141125
R1414 d2 d2 0.1255
R1415 d2 d2 0.063
R1416 d3.n0 d3.t1 556.78
R1417 d3.t1 d3 547.24
R1418 d3 d3.t0 372.113
R1419 d3.n0 d3 9.54008
R1420 d3 d3.n0 0.141125
R1421 d3 d3 0.1255
R1422 d3 d3 0.063
R1423 d4.n0 d4.t1 556.78
R1424 d4.t1 d4 547.24
R1425 d4 d4.t0 372.113
R1426 d4.n0 d4 9.54008
R1427 d4 d4.n0 0.141125
R1428 d4 d4 0.1255
R1429 d4 d4 0.063
R1430 d5.n0 d5.t1 556.78
R1431 d5.t1 d5 547.24
R1432 d5 d5.t0 372.113
R1433 d5.n0 d5 9.54008
R1434 d5 d5.n0 0.141125
R1435 d5 d5 0.1255
R1436 d5 d5 0.063
R1437 d6.n0 d6.t1 556.78
R1438 d6.t1 d6 547.24
R1439 d6 d6.t0 372.113
R1440 d6.n0 d6 9.54008
R1441 d6 d6.n0 0.141125
R1442 d6 d6 0.1255
R1443 d6 d6 0.063
R1444 q0 q0 5.30089
R1445 q0 q0 2.61734
R1446 q1 q1 5.30089
R1447 q1 q1 2.61734
R1448 q2 q2 5.30089
R1449 q2 q2 2.61734
C0 buffer_8/in buffer_1/inv_1/vin 0
C1 tmux_2to1_1/XM5/G tmux_2to1_3/B 0
C2 vdd buffer_5/out 1.92707f
C3 buffer_5/out buffer_4/out 1.95899f
C4 d3 d2 0.00435f
C5 buffer_3/inv_1/vin buffer_4/inv_1/vin 0.00438f
C6 vdd d2 0.07265f
C7 vdd tmux_2to1_3/A 0.31099f
C8 buffer_5/out R1/m1_n100_n100# 0.01185f
C9 R1/R1 buffer_7/in 0.00295f
C10 tmux_2to1_3/A buffer_4/out 0.6033f
C11 buffer_2/inv_1/vin tmux_2to1_3/B 0
C12 buffer_7/in tmux_2to1_3/XM5/G 0.01403f
C13 tmux_2to1_2/XM5/G buffer_5/out 0.09828f
C14 R1/R1 tmux_2to1_3/XM5/G 0
C15 buffer_5/out buffer_6/out 0.48724f
C16 tmux_2to1_0/XM5/G buffer_7/in 0.00597f
C17 vdd buffer_8/inv_1/vin 0.02538f
C18 buffer_5/inv_1/vin buffer_4/inv_1/vin 0.00435f
C19 buffer_8/in buffer_5/out 0.33947f
C20 R1/R1 tmux_2to1_0/XM5/G 0.0674f
C21 buffer_2/out tmux_2to1_3/B 0.04026f
C22 buffer_8/in tmux_2to1_3/A 0.1382f
C23 vdd buffer_3/inv_1/vin 0.32836f
C24 buffer_1/out buffer_1/inv_1/vin 0.0086f
C25 buffer_4/out buffer_3/inv_1/vin 0
C26 buffer_0/out tmux_2to1_3/A 0.05826f
C27 vdd buffer_0/inv_1/vin 0.32203f
C28 R1/m1_n100_n100# buffer_3/inv_1/vin 0.00103f
C29 vdd tmux_2to1_1/XM5/G 0.04059f
C30 buffer_8/in buffer_8/inv_1/vin 0.01384f
C31 buffer_6/out buffer_3/inv_1/vin 0
C32 tmux_2to1_1/XM5/G buffer_4/out 0.02598f
C33 vdd buffer_5/inv_1/vin 0.32846f
C34 R1/R1 R1/R2 0.03366f
C35 tmux_2to1_3/A q0 0
C36 d6 d5 0.00438f
C37 vdd buffer_2/inv_1/vin 0.32649f
C38 tmux_2to1_2/XM5/G tmux_2to1_1/XM5/G 0.00433f
C39 buffer_1/out buffer_5/out 0.05669f
C40 buffer_1/out tmux_2to1_3/A 0
C41 buffer_0/out buffer_0/inv_1/vin 0.00873f
C42 buffer_6/out buffer_5/inv_1/vin 0
C43 buffer_8/in tmux_2to1_1/XM5/G 0.12457f
C44 buffer_9/inv_1/vin buffer_8/inv_1/vin 0.00438f
C45 vdd buffer_2/out 0.64599f
C46 buffer_2/out buffer_4/out 0.0018f
C47 d1 d0 0.00435f
C48 vdd buffer_7/inv_1/vin 0.02382f
C49 buffer_7/inv_1/vin buffer_4/out 0.00238f
C50 tmux_2to1_2/XM5/G buffer_2/out 0.14365f
C51 q1 tmux_2to1_3/B 0
C52 buffer_2/out buffer_6/out 0.01539f
C53 vdd tmux_2to1_3/B 1.44834f
C54 R1/R1 d0 0
C55 buffer_4/out tmux_2to1_3/B 0.27938f
C56 tmux_2to1_1/XM5/G buffer_1/out 0.18587f
C57 buffer_6/inv_1/vin buffer_5/inv_1/vin 0.00438f
C58 tmux_2to1_2/XM5/G tmux_2to1_3/B 0.03416f
C59 tmux_2to1_0/XM5/G d0 0
C60 buffer_6/out tmux_2to1_3/B 0.18281f
C61 q2 tmux_2to1_3/B 0
C62 R1/R1 buffer_1/inv_1/vin 0.02062f
C63 vdd buffer_4/inv_1/vin 0.32846f
C64 buffer_8/in tmux_2to1_3/B 0.28179f
C65 buffer_4/out buffer_4/inv_1/vin 0.00786f
C66 d1 d2 0.00438f
C67 d4 d3 0.00438f
C68 buffer_6/out buffer_4/inv_1/vin 0
C69 vdd q1 0.01294f
C70 buffer_7/in buffer_5/out 0.00264f
C71 vdd d4 0.07265f
C72 d4 buffer_4/out 0.00132f
C73 vdd d3 0.07265f
C74 R1/R1 buffer_5/out 0.55887f
C75 buffer_5/out tmux_2to1_3/XM5/G 0.01262f
C76 buffer_7/in tmux_2to1_3/A 0.38438f
C77 buffer_9/inv_1/vin tmux_2to1_3/B 0.00176f
C78 vdd buffer_4/out 1.75243f
C79 R1/R1 d2 0.00119f
C80 R1/R1 tmux_2to1_3/A 0.0222f
C81 tmux_2to1_3/XM5/G tmux_2to1_3/A 0.04146f
C82 vdd R1/m1_n100_n100# 0.01544f
C83 R1/m1_n100_n100# buffer_4/out 0.00131f
C84 buffer_1/out tmux_2to1_3/B 0
C85 tmux_2to1_2/XM5/G vdd 0.05427f
C86 tmux_2to1_2/XM5/G buffer_4/out 0.07683f
C87 buffer_7/in buffer_8/inv_1/vin 0
C88 buffer_8/in q1 0
C89 vdd buffer_6/out 2.9681f
C90 tmux_2to1_0/XM5/G tmux_2to1_3/A 0.08101f
C91 vdd q2 0.01294f
C92 buffer_6/out buffer_4/out 1.41424f
C93 vdd buffer_8/in 0.52301f
C94 buffer_8/in buffer_4/out 0.18314f
C95 buffer_6/out R1/m1_n100_n100# 0
C96 R1/R1 buffer_3/inv_1/vin 0.00894f
C97 vdd buffer_0/out 0.83616f
C98 tmux_2to1_2/XM5/G buffer_6/out 0.02333f
C99 buffer_0/out buffer_4/out 0.0414f
C100 R1/R1 buffer_0/inv_1/vin 0.01886f
C101 buffer_5/out R1/R2 0.01212f
C102 tmux_2to1_1/XM5/G buffer_7/in 0
C103 vdd q0 0.01294f
C104 R1/R1 tmux_2to1_1/XM5/G 0.13419f
C105 buffer_9/inv_1/vin vdd 0.03021f
C106 tmux_2to1_0/XM5/G buffer_0/inv_1/vin 0
C107 R1/R1 buffer_2/inv_1/vin 0.02182f
C108 vdd buffer_6/inv_1/vin 0.32835f
C109 vdd buffer_1/out 0.83708f
C110 tmux_2to1_0/XM5/G tmux_2to1_1/XM5/G 0.00433f
C111 buffer_1/out buffer_4/out 0.00456f
C112 buffer_9/inv_1/vin buffer_6/out 0.00222f
C113 buffer_6/inv_1/vin buffer_6/out 0.00786f
C114 R1/R1 buffer_2/out 0.2789f
C115 buffer_7/inv_1/vin buffer_7/in 0.00796f
C116 buffer_8/in buffer_1/out 0.06403f
C117 vdd d6 0.07265f
C118 d0 tmux_2to1_3/A 0
C119 buffer_5/out d5 0.00133f
C120 buffer_7/in tmux_2to1_3/B 0.20877f
C121 R1/R1 tmux_2to1_3/B 0.24354f
C122 tmux_2to1_3/XM5/G tmux_2to1_3/B 0.0457f
C123 d6 buffer_6/out 0.00132f
C124 d1 vdd 0.07265f
C125 q1 buffer_7/in 0
C126 buffer_5/out tmux_2to1_3/A 0.00456f
C127 buffer_0/inv_1/vin buffer_1/inv_1/vin 0.00435f
C128 vdd buffer_7/in 0.23539f
C129 R1/R1 d3 0
C130 buffer_7/in buffer_4/out 0.04488f
C131 vdd R1/R1 2.20161f
C132 vdd tmux_2to1_3/XM5/G 0.0495f
C133 R1/R1 buffer_4/out 0.26729f
C134 d1 buffer_8/in 0
C135 tmux_2to1_3/XM5/G buffer_4/out 0.04713f
C136 R1/R1 R1/m1_n100_n100# 0.04565f
C137 buffer_5/out buffer_8/inv_1/vin 0
C138 tmux_2to1_2/XM5/G R1/R1 0.26532f
C139 vdd tmux_2to1_0/XM5/G 0.05854f
C140 buffer_2/inv_1/vin buffer_1/inv_1/vin 0.00438f
C141 buffer_5/out buffer_3/inv_1/vin 0
C142 tmux_2to1_0/XM5/G buffer_4/out 0.02654f
C143 R1/R1 buffer_6/out 0.20693f
C144 R1/R1 q2 0
C145 buffer_8/in buffer_7/in 0.24628f
C146 R1/R1 buffer_8/in 0.07792f
C147 buffer_7/in buffer_0/out 0
C148 buffer_8/in tmux_2to1_3/XM5/G 0.34642f
C149 tmux_2to1_3/A buffer_0/inv_1/vin 0
C150 R1/R1 buffer_0/out 0.11396f
C151 tmux_2to1_1/XM5/G buffer_5/out 0.02579f
C152 buffer_5/out buffer_5/inv_1/vin 0.00827f
C153 vdd R1/R2 0.32828f
C154 d1 buffer_1/out 0.00148f
C155 R1/R2 buffer_4/out 0.00232f
C156 tmux_2to1_1/XM5/G tmux_2to1_3/A 0
C157 buffer_7/in q0 0
C158 tmux_2to1_0/XM5/G buffer_0/out 0.18135f
C159 R1/R2 R1/m1_n100_n100# 0.0386f
C160 buffer_9/inv_1/vin R1/R1 0.00349f
C161 buffer_1/out buffer_7/in 0
C162 buffer_6/out R1/R2 0.00154f
C163 R1/R1 buffer_1/out 0.22519f
C164 buffer_1/out tmux_2to1_3/XM5/G 0
C165 buffer_5/out buffer_2/out 0.05213f
C166 buffer_2/out d2 0
C167 buffer_2/inv_1/vin buffer_3/inv_1/vin 0.00435f
C168 buffer_7/inv_1/vin tmux_2to1_3/A 0
C169 buffer_5/out tmux_2to1_3/B 0.16421f
C170 vdd d0 0.0683f
C171 d4 d5 0.00435f
C172 buffer_7/inv_1/vin buffer_8/inv_1/vin 0.00435f
C173 d2 tmux_2to1_3/B 0
C174 tmux_2to1_3/A tmux_2to1_3/B 0.0101f
C175 vdd d5 0.07265f
C176 vdd buffer_1/inv_1/vin 0.32649f
C177 buffer_5/out buffer_4/inv_1/vin 0
C178 buffer_8/inv_1/vin tmux_2to1_3/B 0.00974f
C179 d0 buffer_0/out 0.0015f
C180 buffer_2/inv_1/vin buffer_2/out 0.00356f
C181 d1 R1/R1 0
C182 vdd.n0 vss 0.03534f
C183 vdd.n1 vss 0.00121f
C184 vdd.n2 vss 0.00532f
C185 vdd.n3 vss 0.00788f
C186 vdd.n4 vss 0.00506f
C187 vdd.n5 vss 0.00788f
C188 vdd.n6 vss 0.05932f
C189 vdd.n7 vss 0.00532f
C190 vdd.n8 vss 0.00506f
C191 vdd.n9 vss 0.00506f
C192 vdd.n10 vss 0.00506f
C193 vdd.n11 vss 0.05932f
C194 vdd.n12 vss 0.00524f
C195 vdd.n13 vss 0.00524f
C196 vdd.n14 vss 0.05932f
C197 vdd.n15 vss 0.00808f
C198 vdd.n16 vss 0.00808f
C199 vdd.n17 vss 0.00282f
C200 vdd.n18 vss 0.00405f
C201 vdd.n19 vss 0.06499f
C202 vdd.n20 vss 0.00808f
C203 vdd.n21 vss 0.00808f
C204 vdd.n22 vss 0.02805f
C205 vdd.n23 vss 0.00627f
C206 vdd.n24 vss 0.03709f
C207 vdd.n25 vss 0.00389f
C208 vdd.n26 vss 0.00405f
C209 vdd.n28 vss 0.05178f
C210 vdd.n29 vss 0.00788f
C211 vdd.n30 vss 0.00788f
C212 vdd.n31 vss 0.00788f
C213 vdd.n32 vss 0.04918f
C214 vdd.n33 vss 0.04918f
C215 vdd.n34 vss 0.00788f
C216 vdd.n35 vss 0.00788f
C217 vdd.n36 vss 0.00788f
C218 vdd.n37 vss 0.00788f
C219 vdd.n38 vss 0.24742f
C220 vdd.n39 vss 0.05932f
C221 vdd.n40 vss 0.24742f
C222 vdd.n41 vss 0.00788f
C223 vdd.n42 vss 0.00788f
C224 vdd.n43 vss 0.00524f
C225 vdd.n44 vss 0.00506f
C226 vdd.n45 vss 0.00532f
C227 vdd.n46 vss 0.00532f
C228 vdd.n47 vss 0.00506f
C229 vdd.n48 vss 0.00241f
C230 vdd.n49 vss 0.05932f
C231 vdd.n50 vss 0.00241f
C232 vdd.n51 vss 0.00506f
C233 vdd.n52 vss 0.00524f
C234 vdd.n53 vss 0.05932f
C235 vdd.n54 vss 0.00808f
C236 vdd.n55 vss 0.00808f
C237 vdd.n56 vss 0.00405f
C238 vdd.n57 vss 0.00282f
C239 vdd.n58 vss 0.06499f
C240 vdd.n59 vss 0.00808f
C241 vdd.n60 vss 0.00808f
C242 vdd.n61 vss 0.00405f
C243 vdd.n62 vss 0.00631f
C244 vdd.n63 vss 0.02805f
C245 vdd.n64 vss 0.02805f
C246 vdd.n65 vss 0.00627f
C247 vdd.n66 vss 0.00282f
C248 vdd.n68 vss 0.05178f
C249 vdd.n69 vss 0.00788f
C250 vdd.n70 vss 0.00788f
C251 vdd.n71 vss 0.00788f
C252 vdd.n72 vss 0.04918f
C253 vdd.n73 vss 0.04918f
C254 vdd.n74 vss 0.00788f
C255 vdd.n75 vss 0.00788f
C256 vdd.n76 vss 0.00788f
C257 vdd.n77 vss 0.00788f
C258 vdd.n78 vss 0.04956f
C259 vdd.n79 vss 0.04956f
C260 vdd.n80 vss 0.05932f
C261 vdd.n81 vss 0.00524f
C262 vdd.n82 vss 0.00524f
C263 vdd.n83 vss 0.00506f
C264 vdd.n84 vss 0.0012f
C265 vdd.n85 vss 0.0176f
C266 vdd.n86 vss 0.12744f
C267 vdd.n87 vss 1.3687f
C268 vdd.n88 vss 0.00282f
C269 vdd.n89 vss 0.0561f
C270 vdd.n90 vss 0.00405f
C271 vdd.n91 vss 0.00808f
C272 vdd.n92 vss 0.00808f
C273 vdd.n93 vss 0.40094f
C274 vdd.n94 vss 0.00788f
C275 vdd.n95 vss 0.40094f
C276 vdd.n96 vss 0.00788f
C277 vdd.n97 vss 0.00788f
C278 vdd.n98 vss 0.00808f
C279 vdd.n99 vss 0.00808f
C280 vdd.n100 vss 0.00788f
C281 vdd.n101 vss 0.00405f
C282 vdd.n102 vss 0.00808f
C283 vdd.n103 vss 0.00808f
C284 vdd.n104 vss 0.40094f
C285 vdd.n105 vss 0.00788f
C286 vdd.n106 vss 0.00788f
C287 vdd.n107 vss 0.00788f
C288 vdd.n108 vss 0.40094f
C289 vdd.n109 vss 0.00808f
C290 vdd.n110 vss 0.00808f
C291 vdd.n111 vss 0.00405f
C292 vdd.n112 vss 0.00788f
C293 vdd.n113 vss 0.00788f
C294 vdd.n114 vss 0.00788f
C295 vdd.n115 vss 0.6218f
C296 vdd.n116 vss 0.00788f
C297 vdd.n117 vss 0.00788f
C298 vdd.n118 vss 0.00282f
C299 vdd.n119 vss 0.0561f
C300 vdd.n120 vss 0.01254f
C301 vdd.n121 vss 0.00282f
C302 vdd.n122 vss 0.00405f
C303 vdd.n123 vss 0.00788f
C304 vdd.n124 vss 0.00788f
C305 vdd.n125 vss 0.6218f
C306 vdd.n126 vss 0.00788f
C307 vdd.n127 vss 0.00788f
C308 vdd.n128 vss 0.00282f
C309 vdd.n129 vss 0.06342f
C310 vdd.n130 vss 0.58772f
C311 vdd.n131 vss 0.00282f
C312 vdd.n132 vss 0.0561f
C313 vdd.n133 vss 0.00405f
C314 vdd.n134 vss 0.00808f
C315 vdd.n135 vss 0.00808f
C316 vdd.n136 vss 0.40094f
C317 vdd.n137 vss 0.00788f
C318 vdd.n138 vss 0.40094f
C319 vdd.n139 vss 0.00788f
C320 vdd.n140 vss 0.00788f
C321 vdd.n141 vss 0.00808f
C322 vdd.n142 vss 0.00808f
C323 vdd.n143 vss 0.00788f
C324 vdd.n144 vss 0.00405f
C325 vdd.n145 vss 0.00808f
C326 vdd.n146 vss 0.00808f
C327 vdd.n147 vss 0.40094f
C328 vdd.n148 vss 0.00788f
C329 vdd.n149 vss 0.00788f
C330 vdd.n150 vss 0.00788f
C331 vdd.n151 vss 0.40094f
C332 vdd.n152 vss 0.00808f
C333 vdd.n153 vss 0.00808f
C334 vdd.n154 vss 0.00405f
C335 vdd.n155 vss 0.00788f
C336 vdd.n156 vss 0.00788f
C337 vdd.n157 vss 0.00788f
C338 vdd.n158 vss 0.6218f
C339 vdd.n159 vss 0.00788f
C340 vdd.n160 vss 0.00788f
C341 vdd.n161 vss 0.00282f
C342 vdd.n162 vss 0.0561f
C343 vdd.n163 vss 0.01254f
C344 vdd.n164 vss 0.00282f
C345 vdd.n165 vss 0.00405f
C346 vdd.n166 vss 0.00788f
C347 vdd.n167 vss 0.00788f
C348 vdd.n168 vss 0.6218f
C349 vdd.n169 vss 0.00788f
C350 vdd.n170 vss 0.00788f
C351 vdd.n171 vss 0.00282f
C352 vdd.n172 vss 0.06073f
C353 vdd.n173 vss 0.31058f
C354 vdd.n174 vss 1.84762f
C355 vdd.n175 vss 0.0012f
C356 vdd.n176 vss 0.07068f
C357 vdd.n177 vss 0.00121f
C358 vdd.n178 vss 0.00532f
C359 vdd.n179 vss 0.00788f
C360 vdd.n180 vss 0.00506f
C361 vdd.n181 vss 0.00788f
C362 vdd.n182 vss 0.11864f
C363 vdd.n183 vss 0.00524f
C364 vdd.n184 vss 0.00788f
C365 vdd.n185 vss 0.11864f
C366 vdd.n186 vss 0.00808f
C367 vdd.n187 vss 0.00808f
C368 vdd.n188 vss 0.00788f
C369 vdd.n189 vss 0.00282f
C370 vdd.n190 vss 0.00282f
C371 vdd.n191 vss 0.0561f
C372 vdd.n192 vss 0.00405f
C373 vdd.n193 vss 0.00808f
C374 vdd.n194 vss 0.00808f
C375 vdd.n195 vss 0.11864f
C376 vdd.n196 vss 0.00808f
C377 vdd.n197 vss 0.00808f
C378 vdd.n198 vss 0.00405f
C379 vdd.n199 vss 0.00808f
C380 vdd.n200 vss 0.00808f
C381 vdd.n201 vss 0.00405f
C382 vdd.n202 vss 0.00788f
C383 vdd.n203 vss 0.00788f
C384 vdd.n204 vss 0.00788f
C385 vdd.n205 vss 0.00788f
C386 vdd.n206 vss 0.09837f
C387 vdd.n207 vss 0.00788f
C388 vdd.n208 vss 0.00788f
C389 vdd.n209 vss 0.09837f
C390 vdd.n210 vss 0.00788f
C391 vdd.n211 vss 0.00788f
C392 vdd.n212 vss 0.00788f
C393 vdd.n213 vss 0.00788f
C394 vdd.n214 vss 0.09912f
C395 vdd.n215 vss 0.00788f
C396 vdd.n216 vss 0.00788f
C397 vdd.n217 vss 0.00282f
C398 vdd.n218 vss 0.01254f
C399 vdd.n219 vss 0.0561f
C400 vdd.n220 vss 0.01262f
C401 vdd.n221 vss 0.00282f
C402 vdd.n222 vss 0.00405f
C403 vdd.n223 vss 0.00788f
C404 vdd.n224 vss 0.00788f
C405 vdd.n225 vss 0.09912f
C406 vdd.n226 vss 0.09912f
C407 vdd.n227 vss 0.00524f
C408 vdd.n228 vss 0.00532f
C409 vdd.n229 vss 0.00506f
C410 vdd.n230 vss 0.00506f
C411 vdd.n231 vss 0.00506f
C412 vdd.n232 vss 0.11864f
C413 vdd.n233 vss 0.00241f
C414 vdd.n234 vss 0.00241f
C415 vdd.n235 vss 0.00506f
C416 vdd.n236 vss 0.00506f
C417 vdd.n237 vss 0.00524f
C418 vdd.n238 vss 0.00506f
C419 vdd.n239 vss 0.00532f
C420 vdd.n240 vss 0.00532f
C421 vdd.n241 vss 0.00506f
C422 vdd.n242 vss 0.00524f
C423 vdd.n243 vss 0.00788f
C424 vdd.n244 vss 0.00788f
C425 vdd.n245 vss 0.00506f
C426 vdd.n246 vss 0.00506f
C427 vdd.n247 vss 0.00788f
C428 vdd.n248 vss 0.00788f
C429 vdd.n249 vss 0.11864f
C430 vdd.n250 vss 0.00524f
C431 vdd.n251 vss 0.00524f
C432 vdd.n252 vss 0.00532f
C433 vdd.n253 vss 0.00121f
C434 vdd.n254 vss 0.00282f
C435 vdd.n255 vss 0.00405f
C436 vdd.n256 vss 0.00808f
C437 vdd.n257 vss 0.00808f
C438 vdd.n258 vss 0.11864f
C439 vdd.n259 vss 0.00808f
C440 vdd.n260 vss 0.00808f
C441 vdd.n261 vss 0.00405f
C442 vdd.n262 vss 0.11864f
C443 vdd.n263 vss 0.00788f
C444 vdd.n264 vss 0.00808f
C445 vdd.n265 vss 0.00808f
C446 vdd.n266 vss 0.00282f
C447 vdd.n267 vss 0.00405f
C448 vdd.n268 vss 0.00808f
C449 vdd.n269 vss 0.00808f
C450 vdd.n270 vss 0.00788f
C451 vdd.n271 vss 0.0561f
C452 vdd.n272 vss 0.02021f
C453 vdd.n273 vss 0.00282f
C454 vdd.n274 vss 0.00405f
C455 vdd.n275 vss 0.00788f
C456 vdd.n276 vss 0.00788f
C457 vdd.n277 vss 0.09912f
C458 vdd.n278 vss 0.00788f
C459 vdd.n279 vss 0.00788f
C460 vdd.n280 vss 0.00788f
C461 vdd.n281 vss 0.00788f
C462 vdd.n282 vss 0.09837f
C463 vdd.n283 vss 0.00788f
C464 vdd.n284 vss 0.00788f
C465 vdd.n285 vss 0.09837f
C466 vdd.n286 vss 0.00788f
C467 vdd.n287 vss 0.00788f
C468 vdd.n288 vss 0.00788f
C469 vdd.n289 vss 0.00788f
C470 vdd.n290 vss 0.11864f
C471 vdd.n291 vss 0.00524f
C472 vdd.n292 vss 0.00524f
C473 vdd.n293 vss 0.00506f
C474 vdd.n294 vss 0.00506f
C475 vdd.n295 vss 0.00506f
C476 vdd.n296 vss 0.00241f
C477 vdd.n297 vss 0.11864f
C478 vdd.n298 vss 0.00506f
C479 vdd.n299 vss 0.00532f
C480 vdd.n300 vss 0.00506f
C481 vdd.n301 vss 0.00506f
C482 vdd.n302 vss 0.00241f
C483 vdd.n303 vss 0.11864f
C484 vdd.n304 vss 0.11864f
C485 vdd.n305 vss 0.00532f
C486 vdd.n306 vss 0.00532f
C487 vdd.n307 vss 0.00506f
C488 vdd.n308 vss 0.00524f
C489 vdd.n309 vss 0.00788f
C490 vdd.n310 vss 0.00788f
C491 vdd.n311 vss 0.09912f
C492 vdd.n312 vss 0.09912f
C493 vdd.n313 vss 0.00788f
C494 vdd.n314 vss 0.00788f
C495 vdd.n315 vss 0.00282f
C496 vdd.n316 vss 0.01254f
C497 vdd.n317 vss 0.0561f
C498 vdd.n318 vss 0.04477f
C499 vdd.n319 vss 0.03545f
C500 vdd.n320 vss 0.0012f
C501 vdd.n321 vss 0.00506f
C502 vdd.n322 vss 0.00524f
C503 vdd.n323 vss 0.00788f
C504 vdd.n324 vss 0.00788f
C505 vdd.n325 vss 0.09912f
C506 vdd.n326 vss 0.09912f
C507 vdd.n327 vss 0.00524f
C508 vdd.n328 vss 0.00524f
C509 vdd.n329 vss 0.00788f
C510 vdd.n330 vss 0.00506f
C511 vdd.n331 vss 0.00532f
C512 vdd.n332 vss 0.00532f
C513 vdd.n333 vss 0.00506f
C514 vdd.n334 vss 0.00524f
C515 vdd.n335 vss 0.00788f
C516 vdd.n336 vss 0.00524f
C517 vdd.n337 vss 0.11864f
C518 vdd.n338 vss 0.00524f
C519 vdd.n339 vss 0.00506f
C520 vdd.n340 vss 0.00532f
C521 vdd.n341 vss 0.00532f
C522 vdd.n342 vss 0.00506f
C523 vdd.n343 vss 0.00121f
C524 vdd.n344 vss 0.00241f
C525 vdd.n345 vss 0.11864f
C526 vdd.n346 vss 0.00241f
C527 vdd.n347 vss 0.00506f
C528 vdd.n348 vss 0.00524f
C529 vdd.n349 vss 0.11864f
C530 vdd.n350 vss 0.00524f
C531 vdd.n351 vss 0.00524f
C532 vdd.n352 vss 0.00506f
C533 vdd.n353 vss 0.0012f
C534 vdd.n354 vss 0.03534f
C535 vdd.n355 vss 0.01892f
C536 vdd.n356 vss 0.25756f
C537 vdd.n357 vss 0.39762f
C538 tmux_2to1_3/A vss 0.7137f
C539 tmux_2to1_0/XM5/G vss 0.55203f
C540 buffer_9/inv_1/vin vss 0.83718f
C541 q2 vss 0.40182f
C542 buffer_8/inv_1/vin vss 0.83586f
C543 q1 vss 0.40182f
C544 buffer_7/inv_1/vin vss 0.83588f
C545 q0 vss 0.40182f
C546 buffer_6/inv_1/vin vss 0.54713f
C547 buffer_6/out vss 1.02817f
C548 d6 vss 0.42023f
C549 buffer_5/inv_1/vin vss 0.54811f
C550 buffer_5/out vss 1.10288f
C551 d5 vss 0.41693f
C552 vdd vss 82.618f
C553 buffer_4/inv_1/vin vss 0.54811f
C554 buffer_4/out vss 1.13783f
C555 d4 vss 0.41693f
C556 buffer_3/inv_1/vin vss 0.54811f
C557 R1/R2 vss 0.24595f
C558 d3 vss 0.41694f
C559 buffer_2/inv_1/vin vss 0.55981f
C560 buffer_2/out vss 0.38944f
C561 d2 vss 0.41693f
C562 buffer_1/inv_1/vin vss 0.55981f
C563 buffer_1/out vss 0.403f
C564 d1 vss 0.41693f
C565 buffer_0/inv_1/vin vss 0.55981f
C566 buffer_0/out vss 0.40723f
C567 d0 vss 0.42457f
C568 R1/m1_n100_n100# vss 0.11104f
C569 buffer_8/in vss 1.94693f
C570 buffer_7/in vss 1.30882f
C571 tmux_2to1_3/XM5/G vss 0.55181f
C572 R1/R1 vss 4.97016f
C573 tmux_2to1_3/B vss 1.00035f
C574 tmux_2to1_2/XM5/G vss 0.54992f
C575 tmux_2to1_1/XM5/G vss 0.55178f
.ends

