* NGSPICE file created from tt_um_tinyflash_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9 B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_1p41 l=7
C0 R2 R1 0.01325f
C1 R2 B 0.82332f
C2 R1 B 0.82332f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ELBHUY B D S G
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 G D 0.11229f
C1 S D 0.27388f
C2 S G 0.11229f
C3 S B 0.59197f
C4 D B 0.59197f
C5 G B 0.75059f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_VTBKAA B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 S G 0.21915f
C1 S B 0.634f
C2 D S 0.54671f
C3 B G 0.43443f
C4 D G 0.21915f
C5 D B 0.634f
C6 S VSUBS 0.51455f
C7 D VSUBS 0.51455f
C8 G VSUBS 0.36418f
C9 B VSUBS 5.72384f
.ends

.subckt vbias_generation bias_n vdd XR_bias_2/R2 XR_bias_4/R1 XR_bias_3/R2 bias_p
+ vss
XXR_bias_1 vss XR_bias_2/R2 bias_p sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_2 vss XR_bias_3/R2 XR_bias_2/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_3 vss XR_bias_4/R1 XR_bias_3/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_4 vss XR_bias_4/R1 bias_n sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXMn_bias vss bias_n vss bias_n sky130_fd_pr__nfet_01v8_lvt_ELBHUY
XXMp_bias vdd bias_p vdd bias_p vss sky130_fd_pr__pfet_01v8_lvt_VTBKAA
C0 XR_bias_4/R1 XR_bias_3/R2 0
C1 XR_bias_2/R2 bias_p 0.05112f
C2 XR_bias_2/R2 vdd 0.01866f
C3 vdd bias_p 0.22745f
C4 XR_bias_2/R2 XR_bias_4/R1 0.06887f
C5 XR_bias_2/R2 XR_bias_3/R2 0
C6 XR_bias_4/R1 bias_p 0
C7 bias_p XR_bias_3/R2 0.06932f
C8 XR_bias_4/R1 bias_n 0
C9 bias_n XR_bias_3/R2 0.06908f
C10 vdd vss 6.78775f
C11 bias_n vss 2.48381f
C12 XR_bias_4/R1 vss 1.63605f
C13 XR_bias_3/R2 vss 1.57785f
C14 XR_bias_2/R2 vss 1.57097f
C15 bias_p vss 1.64123f
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_JT48NU B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_5p73 l=5.73
C0 R2 R1 0.06813f
C1 R2 B 1.74197f
C2 R1 B 1.74197f
.ends

.subckt res_ladder_vref ref2 ref5 ref6 vref ref3 ref1 ref0 ref4 vss
XXR1 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR2 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR10 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR3 vss ref6 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR4 vss ref4 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR5 vss ref4 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR6 vss ref2 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR7 vss ref2 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR8 vss ref0 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR9 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
C0 ref6 ref5 0
C1 ref2 ref4 0.06887f
C2 ref3 ref4 0
C3 ref6 ref4 0.06887f
C4 ref2 ref3 0
C5 ref2 ref0 0.06887f
C6 ref5 ref4 0
C7 vref ref6 0.16095f
C8 ref2 ref1 0
C9 vref ref5 0.06887f
C10 ref3 ref1 0.06887f
C11 ref3 ref5 0.06887f
C12 ref1 ref0 0
C13 ref1 vss 3.4889f
C14 ref2 vss 3.42003f
C15 ref3 vss 3.42003f
C16 ref4 vss 3.42003f
C17 ref5 vss 3.42003f
C18 ref6 vss 5.161f
C19 ref0 vss 5.32418f
C20 vref vss 4.57377f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MMMA4V a_n260_n698# a_100_n500# a_n158_n500# a_n100_n588#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n698# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 a_n158_n500# a_n100_n588# 0.11229f
C1 a_n158_n500# a_100_n500# 0.27388f
C2 a_n100_n588# a_100_n500# 0.11229f
C3 a_100_n500# a_n260_n698# 0.5905f
C4 a_n158_n500# a_n260_n698# 0.5905f
C5 a_n100_n588# a_n260_n698# 0.7183f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_5VNMZ8 a_n100_n897# a_100_n800# w_n296_n1019#
+ a_n158_n800# VSUBS
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n296_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
C0 a_n100_n897# w_n296_n1019# 0.43443f
C1 a_n100_n897# a_n158_n800# 0.17641f
C2 a_100_n800# a_n100_n897# 0.17641f
C3 w_n296_n1019# a_n158_n800# 0.51205f
C4 a_100_n800# w_n296_n1019# 0.51205f
C5 a_100_n800# a_n158_n800# 0.43758f
C6 a_100_n800# VSUBS 0.41369f
C7 a_n158_n800# VSUBS 0.41369f
C8 a_n100_n897# VSUBS 0.36418f
C9 w_n296_n1019# VSUBS 4.82082f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHMAL2 a_n260_n574# a_100_n400# a_n158_n400# a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n260_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
C0 a_n158_n400# a_n100_n488# 0.09092f
C1 a_n158_n400# a_100_n400# 0.21931f
C2 a_n100_n488# a_100_n400# 0.09092f
C3 a_100_n400# a_n260_n574# 0.48057f
C4 a_n158_n400# a_n260_n574# 0.48057f
C5 a_n100_n488# a_n260_n574# 0.74751f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GUWLND a_n158_n1000# a_n100_n1097# w_n296_n1219#
+ a_100_n1000# VSUBS
X0 a_100_n1000# a_n100_n1097# a_n158_n1000# w_n296_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 a_n100_n1097# w_n296_n1219# 0.43443f
C1 a_n100_n1097# a_n158_n1000# 0.21915f
C2 a_100_n1000# a_n100_n1097# 0.21915f
C3 w_n296_n1219# a_n158_n1000# 0.634f
C4 a_100_n1000# w_n296_n1219# 0.634f
C5 a_100_n1000# a_n158_n1000# 0.54671f
C6 a_100_n1000# VSUBS 0.51455f
C7 a_n158_n1000# VSUBS 0.51455f
C8 a_n100_n1097# VSUBS 0.36418f
C9 w_n296_n1219# VSUBS 5.72384f
.ends

.subckt comp_p vinp vinn vbias_p vdd tail vout latch_right out_left latch_left vss
XXMn_cs_left vss latch_right vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_out out_left vdd vdd vout vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_diode_left1 vss latch_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_AHMAL2
XXMn_cs_right1 vss latch_left vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_diode_right vss latch_right vss latch_right sky130_fd_pr__nfet_01v8_lvt_AHMAL2
Xsky130_fd_pr__pfet_01v8_lvt_5VNMZ8_0 out_left vdd vdd out_left vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_out_left vss out_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_out_right vss vout vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_tail tail vbias_p vdd vdd vss sky130_fd_pr__pfet_01v8_lvt_GUWLND
X0 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X1 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X2 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X3 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X4 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X5 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X6 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X7 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
C0 vout vinp 0.03655f
C1 vinn latch_right 3.53507f
C2 out_left vdd 2.99708f
C3 latch_left vdd 1.3971f
C4 vbias_p vout 0.14426f
C5 out_left vinp 0.22514f
C6 vdd vinn 2.30474f
C7 latch_left vinp 0.5043f
C8 vbias_p out_left 0.84152f
C9 vbias_p latch_left 0.00103f
C10 vinn vinp 1.25697f
C11 tail latch_right 8.8942f
C12 vbias_p vinn 0.00222f
C13 vdd tail 2.22915f
C14 out_left vout 0.6058f
C15 latch_left vout 0.14014f
C16 tail vinp 2.91757f
C17 vdd latch_right 1.44611f
C18 vout vinn 0.12978f
C19 out_left latch_left 0.73463f
C20 vbias_p tail 0.65167f
C21 latch_right vinp 0.51311f
C22 out_left vinn 0.08183f
C23 latch_left vinn 1.33911f
C24 vbias_p latch_right 0.00109f
C25 vdd vinp 4.26352f
C26 vout tail 0.00803f
C27 vbias_p vdd 2.11961f
C28 vout latch_right 0.72835f
C29 out_left tail 0.00652f
C30 vbias_p vinp 0.03011f
C31 latch_left tail 8.82993f
C32 out_left latch_right 0.1431f
C33 vout vdd 1.62919f
C34 vinn tail 0.82695f
C35 latch_left latch_right 5.15792f
C36 vinp vss 0.4258f
C37 vinn vss 0.50566f
C38 tail vss 1.09774f
C39 vbias_p vss 0.82905f
C40 vdd vss 43.54159f
C41 vout vss 3.2381f
C42 latch_right vss 4.74799f
C43 out_left vss 3.38408f
C44 latch_left vss 5.11722f
.ends

.subckt sky130_fd_pr__pfet_01v8_A6MZLZ B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 S G 0.02934f
C1 S D 0.32105f
C2 S B 0.14266f
C3 G D 0.02934f
C4 G B 0.24043f
C5 D B 0.14266f
C6 S VSUBS 0.09023f
C7 D VSUBS 0.09023f
C8 G VSUBS 0.11914f
C9 B VSUBS 1.5811f
.ends

.subckt sky130_fd_pr__nfet_01v8_MH3LLV B D S G
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 D S 0.16211f
C1 D G 0.02545f
C2 S G 0.02545f
C3 S B 0.1317f
C4 D B 0.1317f
C5 G B 0.34289f
.ends

.subckt tmux_2to1 Y vdd XM5/G A B S vss
XXM1 vdd vdd XM5/G S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM2 vss vss XM5/G S sky130_fd_pr__nfet_01v8_MH3LLV
XXM3 vdd A Y S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM4 vss A Y XM5/G sky130_fd_pr__nfet_01v8_MH3LLV
XXM5 vdd Y B XM5/G vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM6 vss Y B S sky130_fd_pr__nfet_01v8_MH3LLV
C0 vdd XM5/G 0.17343f
C1 XM5/G A 0.66126f
C2 XM5/G S 0.4752f
C3 B XM5/G 0.09611f
C4 vdd A 0.05809f
C5 vdd S 0.27839f
C6 XM5/G Y 0.31571f
C7 vdd B 0.11322f
C8 A S 0.09932f
C9 vdd Y 0.18933f
C10 B S 0.0426f
C11 A Y 0.03022f
C12 S Y 0.13093f
C13 B Y 0.03022f
C14 B vss 0.39578f
C15 S vss 1.22376f
C16 Y vss 0.38976f
C17 XM5/G vss 0.68597f
C18 vdd vss 4.09633f
C19 A vss 0.18036f
.ends

.subckt sky130_fd_pr__res_generic_m1_SPQYYJ R1 R2 m1_n100_n100# VSUBS
R0 R1 R2 sky130_fd_pr__res_generic_m1 w=1 l=1
C0 R2 VSUBS 0.07104f
C1 R1 VSUBS 0.07104f
C2 m1_n100_n100# VSUBS 0.10692f
.ends

.subckt inv vin vdd vout vss
XXMn vss vss vout vin sky130_fd_pr__nfet_01v8_MH3LLV
XXMp vdd vdd vout vin vss sky130_fd_pr__pfet_01v8_A6MZLZ
C0 vdd vin 0.13776f
C1 vout vin 0.12658f
C2 vdd vout 0.11998f
C3 vin vss 0.56678f
C4 vout vss 0.40687f
C5 vdd vss 1.84972f
.ends

.subckt buffer in out vdd inv_1/vin vss
Xinv_0 in vdd inv_1/vin vss inv
Xinv_1 inv_1/vin vdd out vss inv
C0 in inv_1/vin 0.01628f
C1 in vdd 0.01965f
C2 out inv_1/vin 0.0071f
C3 out vdd 0.00589f
C4 vdd inv_1/vin 0.16476f
C5 inv_1/vin vss 0.60193f
C6 out vss 0.3255f
C7 in vss 0.41789f
C8 vdd vss 3.06334f
.ends

.subckt tmux_7therm_to_3bin d0 d1 d2 d3 d4 d5 d6 q0 q1 q2 buffer_7/inv_1/vin buffer_3/inv_1/vin
+ buffer_2/out buffer_8/inv_1/vin buffer_4/inv_1/vin buffer_0/inv_1/vin buffer_6/out
+ R1/R2 buffer_9/inv_1/vin buffer_0/out buffer_5/inv_1/vin buffer_5/out buffer_1/inv_1/vin
+ tmux_2to1_0/XM5/G tmux_2to1_3/B tmux_2to1_1/XM5/G tmux_2to1_3/A tmux_2to1_2/XM5/G
+ tmux_2to1_3/XM5/G R1/R1 buffer_6/inv_1/vin buffer_2/inv_1/vin R1/m1_n100_n100# buffer_1/out
+ buffer_8/in vdd vss buffer_7/in buffer_4/out
Xtmux_2to1_1 buffer_8/in vdd tmux_2to1_1/XM5/G buffer_1/out buffer_5/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_2 tmux_2to1_3/B vdd tmux_2to1_2/XM5/G buffer_2/out buffer_6/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_3 buffer_7/in vdd tmux_2to1_3/XM5/G tmux_2to1_3/A tmux_2to1_3/B buffer_8/in
+ vss tmux_2to1
XR1 R1/R1 R1/R2 R1/m1_n100_n100# vss sky130_fd_pr__res_generic_m1_SPQYYJ
Xbuffer_0 d0 buffer_0/out vdd buffer_0/inv_1/vin vss buffer
Xbuffer_1 d1 buffer_1/out vdd buffer_1/inv_1/vin vss buffer
Xbuffer_2 d2 buffer_2/out vdd buffer_2/inv_1/vin vss buffer
Xbuffer_3 d3 R1/R2 vdd buffer_3/inv_1/vin vss buffer
Xbuffer_4 d4 buffer_4/out vdd buffer_4/inv_1/vin vss buffer
Xbuffer_5 d5 buffer_5/out vdd buffer_5/inv_1/vin vss buffer
Xbuffer_6 d6 buffer_6/out vdd buffer_6/inv_1/vin vss buffer
Xbuffer_7 buffer_7/in q0 vdd buffer_7/inv_1/vin vss buffer
Xbuffer_8 buffer_8/in q1 vdd buffer_8/inv_1/vin vss buffer
Xbuffer_9 R1/R1 q2 vdd buffer_9/inv_1/vin vss buffer
Xtmux_2to1_0 tmux_2to1_3/A vdd tmux_2to1_0/XM5/G buffer_0/out buffer_4/out R1/R1 vss
+ tmux_2to1
C0 buffer_0/out buffer_7/in 0
C1 vdd tmux_2to1_3/A 0.31099f
C2 buffer_8/inv_1/vin buffer_7/inv_1/vin 0.00435f
C3 R1/R1 tmux_2to1_3/A 0.0222f
C4 vdd buffer_2/inv_1/vin 0.32649f
C5 buffer_6/out tmux_2to1_2/XM5/G 0.02333f
C6 tmux_2to1_3/B q2 0
C7 buffer_5/out buffer_8/inv_1/vin 0
C8 R1/R1 buffer_2/inv_1/vin 0.02182f
C9 d4 d5 0.00435f
C10 tmux_2to1_3/B buffer_4/out 0.27941f
C11 tmux_2to1_3/B tmux_2to1_3/XM5/G 0.0457f
C12 buffer_5/inv_1/vin vdd 0.32846f
C13 tmux_2to1_3/B d2 0
C14 buffer_0/inv_1/vin vdd 0.32203f
C15 buffer_0/inv_1/vin R1/R1 0.01886f
C16 buffer_4/out buffer_7/inv_1/vin 0.00238f
C17 tmux_2to1_3/B buffer_1/out 0
C18 vdd buffer_9/inv_1/vin 0.03021f
C19 buffer_4/inv_1/vin vdd 0.32846f
C20 buffer_5/out buffer_4/out 1.96436f
C21 R1/R1 buffer_9/inv_1/vin 0.00349f
C22 tmux_2to1_3/B buffer_6/out 0.18281f
C23 d3 d2 0.00435f
C24 buffer_5/out tmux_2to1_3/XM5/G 0.01262f
C25 buffer_4/out tmux_2to1_0/XM5/G 0.02654f
C26 d0 tmux_2to1_0/XM5/G 0
C27 buffer_2/out buffer_4/out 0.0018f
C28 d6 vdd 0.07265f
C29 buffer_4/out tmux_2to1_1/XM5/G 0.02598f
C30 buffer_1/out buffer_5/out 0.05669f
C31 buffer_6/out buffer_5/out 0.48773f
C32 R1/R1 vdd 2.2016f
C33 buffer_2/out d2 0
C34 buffer_8/in buffer_7/in 0.24628f
C35 buffer_1/inv_1/vin buffer_8/in 0
C36 buffer_1/out tmux_2to1_1/XM5/G 0.18587f
C37 buffer_4/out tmux_2to1_3/A 0.60354f
C38 buffer_2/out buffer_6/out 0.01539f
C39 buffer_5/out d5 0.00133f
C40 d1 vdd 0.07265f
C41 buffer_8/inv_1/vin buffer_9/inv_1/vin 0.00438f
C42 tmux_2to1_3/XM5/G tmux_2to1_3/A 0.04146f
C43 d0 tmux_2to1_3/A 0
C44 d1 R1/R1 0
C45 buffer_0/out tmux_2to1_0/XM5/G 0.18135f
C46 buffer_3/inv_1/vin buffer_5/out 0
C47 buffer_1/out tmux_2to1_3/A 0
C48 buffer_5/out R1/m1_n100_n100# 0.01185f
C49 q0 tmux_2to1_3/A 0
C50 buffer_4/out buffer_4/inv_1/vin 0.0079f
C51 buffer_8/inv_1/vin vdd 0.02538f
C52 q1 buffer_8/in 0
C53 tmux_2to1_3/B buffer_8/in 0.28179f
C54 buffer_0/out tmux_2to1_3/A 0.05826f
C55 buffer_6/out buffer_5/inv_1/vin 0
C56 R1/R2 buffer_5/out 0.01212f
C57 q2 vdd 0.01294f
C58 q2 R1/R1 0
C59 buffer_6/out buffer_9/inv_1/vin 0.00222f
C60 buffer_6/out buffer_4/inv_1/vin 0
C61 buffer_4/out vdd 1.78677f
C62 q1 buffer_7/in 0
C63 tmux_2to1_3/B buffer_7/in 0.20877f
C64 buffer_4/out R1/R1 0.26729f
C65 buffer_6/inv_1/vin buffer_5/inv_1/vin 0.00438f
C66 tmux_2to1_3/XM5/G vdd 0.0495f
C67 buffer_3/inv_1/vin buffer_2/inv_1/vin 0.00435f
C68 d0 vdd 0.0683f
C69 tmux_2to1_3/XM5/G R1/R1 0
C70 d0 R1/R1 0
C71 buffer_5/out buffer_8/in 0.33947f
C72 buffer_0/inv_1/vin buffer_0/out 0.00873f
C73 d2 vdd 0.07265f
C74 d2 R1/R1 0.00119f
C75 buffer_6/out d6 0.00132f
C76 buffer_7/in buffer_7/inv_1/vin 0.00796f
C77 buffer_1/out vdd 0.83708f
C78 buffer_1/out R1/R1 0.22519f
C79 buffer_5/out buffer_7/in 0.00264f
C80 buffer_6/out vdd 3.00774f
C81 d3 d4 0.00438f
C82 d1 d0 0.00435f
C83 buffer_6/out R1/R1 0.20693f
C84 tmux_2to1_3/B tmux_2to1_2/XM5/G 0.03416f
C85 buffer_8/in tmux_2to1_1/XM5/G 0.12457f
C86 q0 vdd 0.01294f
C87 buffer_7/in tmux_2to1_0/XM5/G 0.00597f
C88 d1 d2 0.00438f
C89 buffer_3/inv_1/vin buffer_4/inv_1/vin 0.00438f
C90 d5 d6 0.00438f
C91 buffer_6/inv_1/vin vdd 0.32835f
C92 d1 buffer_1/out 0.00148f
C93 tmux_2to1_1/XM5/G buffer_7/in 0
C94 d5 vdd 0.07265f
C95 buffer_0/out vdd 0.83616f
C96 buffer_0/out R1/R1 0.11396f
C97 buffer_8/in tmux_2to1_3/A 0.1382f
C98 buffer_5/out tmux_2to1_2/XM5/G 0.09828f
C99 q1 tmux_2to1_3/B 0
C100 buffer_3/inv_1/vin vdd 0.32836f
C101 buffer_3/inv_1/vin R1/R1 0.00894f
C102 buffer_7/in tmux_2to1_3/A 0.38438f
C103 R1/m1_n100_n100# vdd 0.01544f
C104 buffer_2/out tmux_2to1_2/XM5/G 0.14365f
C105 R1/R1 R1/m1_n100_n100# 0.04565f
C106 tmux_2to1_1/XM5/G tmux_2to1_2/XM5/G 0.00433f
C107 buffer_4/out tmux_2to1_3/XM5/G 0.04713f
C108 buffer_1/inv_1/vin buffer_2/inv_1/vin 0.00438f
C109 tmux_2to1_3/B buffer_5/out 0.16421f
C110 R1/R2 vdd 0.32828f
C111 R1/R2 R1/R1 0.03366f
C112 buffer_1/out buffer_4/out 0.00456f
C113 buffer_1/inv_1/vin buffer_0/inv_1/vin 0.00435f
C114 buffer_2/out tmux_2to1_3/B 0.04026f
C115 buffer_6/out buffer_4/out 1.41966f
C116 buffer_1/out tmux_2to1_3/XM5/G 0
C117 tmux_2to1_3/B tmux_2to1_1/XM5/G 0
C118 buffer_8/in vdd 0.52301f
C119 buffer_8/in R1/R1 0.07792f
C120 buffer_4/out buffer_0/out 0.0414f
C121 buffer_2/out buffer_5/out 0.05213f
C122 tmux_2to1_3/B tmux_2to1_3/A 0.0101f
C123 buffer_5/out tmux_2to1_1/XM5/G 0.02579f
C124 buffer_7/in vdd 0.23539f
C125 R1/R1 buffer_7/in 0.00295f
C126 d0 buffer_0/out 0.0015f
C127 tmux_2to1_3/B buffer_2/inv_1/vin 0
C128 d1 buffer_8/in 0
C129 tmux_2to1_1/XM5/G tmux_2to1_0/XM5/G 0.00433f
C130 buffer_1/inv_1/vin vdd 0.32649f
C131 d4 vdd 0.07265f
C132 buffer_3/inv_1/vin buffer_4/out 0
C133 buffer_1/inv_1/vin R1/R1 0.02062f
C134 tmux_2to1_3/A buffer_7/inv_1/vin 0
C135 buffer_6/out buffer_6/inv_1/vin 0.00786f
C136 buffer_4/out R1/m1_n100_n100# 0.00131f
C137 buffer_5/out tmux_2to1_3/A 0.00456f
C138 tmux_2to1_0/XM5/G tmux_2to1_3/A 0.08101f
C139 tmux_2to1_2/XM5/G vdd 0.05427f
C140 tmux_2to1_2/XM5/G R1/R1 0.26532f
C141 tmux_2to1_3/B buffer_9/inv_1/vin 0.00176f
C142 buffer_8/in buffer_8/inv_1/vin 0.01384f
C143 buffer_6/out buffer_3/inv_1/vin 0
C144 tmux_2to1_1/XM5/G tmux_2to1_3/A 0
C145 R1/R2 buffer_4/out 0.00232f
C146 buffer_5/out buffer_5/inv_1/vin 0.00827f
C147 buffer_6/out R1/m1_n100_n100# 0
C148 buffer_2/out buffer_2/inv_1/vin 0.00356f
C149 buffer_8/inv_1/vin buffer_7/in 0
C150 buffer_0/inv_1/vin tmux_2to1_0/XM5/G 0
C151 buffer_5/out buffer_4/inv_1/vin 0
C152 q1 vdd 0.01294f
C153 tmux_2to1_3/B vdd 1.44834f
C154 tmux_2to1_3/B R1/R1 0.24354f
C155 buffer_4/out buffer_8/in 0.18314f
C156 buffer_8/in tmux_2to1_3/XM5/G 0.34642f
C157 buffer_6/out R1/R2 0.00154f
C158 d3 vdd 0.07265f
C159 vdd buffer_7/inv_1/vin 0.02382f
C160 buffer_4/out buffer_7/in 0.04488f
C161 d3 R1/R1 0
C162 buffer_3/inv_1/vin R1/m1_n100_n100# 0.00103f
C163 tmux_2to1_3/XM5/G buffer_7/in 0.01403f
C164 buffer_5/out vdd 1.96257f
C165 buffer_1/out buffer_8/in 0.06403f
C166 buffer_5/out R1/R1 0.55887f
C167 d4 buffer_4/out 0.00133f
C168 buffer_0/inv_1/vin tmux_2to1_3/A 0
C169 vdd tmux_2to1_0/XM5/G 0.05854f
C170 R1/R1 tmux_2to1_0/XM5/G 0.0674f
C171 buffer_1/out buffer_7/in 0
C172 buffer_2/out vdd 0.64599f
C173 buffer_2/out R1/R1 0.2789f
C174 tmux_2to1_1/XM5/G vdd 0.04059f
C175 buffer_4/out tmux_2to1_2/XM5/G 0.07683f
C176 tmux_2to1_1/XM5/G R1/R1 0.13419f
C177 buffer_1/inv_1/vin buffer_1/out 0.0086f
C178 q0 buffer_7/in 0
C179 tmux_2to1_3/B buffer_8/inv_1/vin 0.00974f
C180 R1/R2 R1/m1_n100_n100# 0.0386f
C181 buffer_5/inv_1/vin buffer_4/inv_1/vin 0.00435f
C182 tmux_2to1_3/A vss 0.7137f
C183 tmux_2to1_0/XM5/G vss 0.55203f
C184 buffer_9/inv_1/vin vss 0.83718f
C185 q2 vss 0.40182f
C186 buffer_8/inv_1/vin vss 0.83586f
C187 q1 vss 0.40182f
C188 buffer_7/inv_1/vin vss 0.83588f
C189 q0 vss 0.40182f
C190 buffer_6/inv_1/vin vss 0.54713f
C191 buffer_6/out vss 1.08087f
C192 d6 vss 0.42023f
C193 buffer_5/inv_1/vin vss 0.54811f
C194 buffer_5/out vss 1.1426f
C195 d5 vss 0.41693f
C196 vdd vss 81.61826f
C197 buffer_4/inv_1/vin vss 0.54811f
C198 buffer_4/out vss 1.13891f
C199 d4 vss 0.41693f
C200 buffer_3/inv_1/vin vss 0.54811f
C201 R1/R2 vss 0.24595f
C202 d3 vss 0.41694f
C203 buffer_2/inv_1/vin vss 0.55981f
C204 buffer_2/out vss 0.38944f
C205 d2 vss 0.41693f
C206 buffer_1/inv_1/vin vss 0.55981f
C207 buffer_1/out vss 0.403f
C208 d1 vss 0.41693f
C209 buffer_0/inv_1/vin vss 0.55981f
C210 buffer_0/out vss 0.40723f
C211 d0 vss 0.42457f
C212 R1/m1_n100_n100# vss 0.11104f
C213 buffer_8/in vss 1.94693f
C214 buffer_7/in vss 1.30882f
C215 tmux_2to1_3/XM5/G vss 0.55181f
C216 R1/R1 vss 4.97016f
C217 tmux_2to1_3/B vss 1.00035f
C218 tmux_2to1_2/XM5/G vss 0.54992f
C219 tmux_2to1_1/XM5/G vss 0.55178f
.ends

.subckt flashADC_3bit dout0 dout1 dout2 tmux_7therm_to_3bin_0/buffer_1/out vbias_generation_0/bias_n
+ tmux_7therm_to_3bin_0/buffer_6/inv_1/vin tmux_7therm_to_3bin_0/buffer_2/inv_1/vin
+ comp_p_3/latch_left comp_p_5/tail tmux_7therm_to_3bin_0/buffer_8/in comp_p_2/tail
+ comp_p_4/latch_left tmux_7therm_to_3bin_0/buffer_7/in comp_p_5/latch_left vbias_generation_0/XR_bias_2/R2
+ tmux_7therm_to_3bin_0/R1/m1_n100_n100# tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_2/out tmux_7therm_to_3bin_0/buffer_3/inv_1/vin comp_p_6/latch_left
+ comp_p_1/out_left comp_p_6/tail comp_p_0/latch_right comp_p_1/latch_right comp_p_2/latch_right
+ comp_p_3/latch_right comp_p_3/tail comp_p_4/latch_right comp_p_5/latch_right tmux_7therm_to_3bin_0/buffer_8/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_6/out comp_p_4/out_left comp_p_4/vinn comp_p_6/latch_right
+ comp_p_0/tail tmux_7therm_to_3bin_0/buffer_4/inv_1/vin tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ tmux_7therm_to_3bin_0/R1/R2 comp_p_2/latch_left vbias_generation_0/XR_bias_4/R1
+ tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G d1 comp_p_3/vinn tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G
+ comp_p_2/out_left tmux_7therm_to_3bin_0/buffer_0/out comp_p_0/out_left tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G
+ tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G comp_p_6/vinn tmux_7therm_to_3bin_0/buffer_5/out
+ d2 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin comp_p_4/tail tmux_7therm_to_3bin_0/R1/R1
+ comp_p_0/latch_left tmux_7therm_to_3bin_0/buffer_5/inv_1/vin tmux_7therm_to_3bin_0/buffer_1/inv_1/vin
+ d4 comp_p_5/vinn tmux_7therm_to_3bin_0/tmux_2to1_3/B comp_p_1/tail comp_p_0/vinn
+ vin comp_p_6/out_left tmux_7therm_to_3bin_0/tmux_2to1_3/A comp_p_1/latch_left vdd
+ tmux_7therm_to_3bin_0/buffer_4/out d5 d3 d0 comp_p_1/vinn comp_p_2/vinn vref comp_p_5/out_left
+ vbias_generation_0/XR_bias_3/R2 d6 vss comp_p_3/out_left comp_p_6/vbias_p
Xvbias_generation_0 vbias_generation_0/bias_n vdd vbias_generation_0/XR_bias_2/R2
+ vbias_generation_0/XR_bias_4/R1 vbias_generation_0/XR_bias_3/R2 comp_p_6/vbias_p
+ vss vbias_generation
Xres_ladder_vref_0 comp_p_2/vinn comp_p_5/vinn comp_p_6/vinn vref comp_p_3/vinn comp_p_0/vinn
+ comp_p_1/vinn comp_p_4/vinn vss res_ladder_vref
Xcomp_p_1 vin comp_p_1/vinn comp_p_6/vbias_p vdd comp_p_1/tail d0 comp_p_1/latch_right
+ comp_p_1/out_left comp_p_1/latch_left vss comp_p
Xcomp_p_0 vin comp_p_0/vinn comp_p_6/vbias_p vdd comp_p_0/tail d1 comp_p_0/latch_right
+ comp_p_0/out_left comp_p_0/latch_left vss comp_p
Xcomp_p_2 vin comp_p_2/vinn comp_p_6/vbias_p vdd comp_p_2/tail d2 comp_p_2/latch_right
+ comp_p_2/out_left comp_p_2/latch_left vss comp_p
Xcomp_p_3 vin comp_p_3/vinn comp_p_6/vbias_p vdd comp_p_3/tail d3 comp_p_3/latch_right
+ comp_p_3/out_left comp_p_3/latch_left vss comp_p
Xcomp_p_4 vin comp_p_4/vinn comp_p_6/vbias_p vdd comp_p_4/tail d4 comp_p_4/latch_right
+ comp_p_4/out_left comp_p_4/latch_left vss comp_p
Xcomp_p_5 vin comp_p_5/vinn comp_p_6/vbias_p vdd comp_p_5/tail d5 comp_p_5/latch_right
+ comp_p_5/out_left comp_p_5/latch_left vss comp_p
Xcomp_p_6 vin comp_p_6/vinn comp_p_6/vbias_p vdd comp_p_6/tail d6 comp_p_6/latch_right
+ comp_p_6/out_left comp_p_6/latch_left vss comp_p
Xtmux_7therm_to_3bin_0 d0 d1 d2 d3 d4 d5 d6 dout0 dout1 dout2 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_3/inv_1/vin tmux_7therm_to_3bin_0/buffer_2/out tmux_7therm_to_3bin_0/buffer_8/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_4/inv_1/vin tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_6/out tmux_7therm_to_3bin_0/R1/R2 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_0/out tmux_7therm_to_3bin_0/buffer_5/inv_1/vin tmux_7therm_to_3bin_0/buffer_5/out
+ tmux_7therm_to_3bin_0/buffer_1/inv_1/vin tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G
+ tmux_7therm_to_3bin_0/tmux_2to1_3/B tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G tmux_7therm_to_3bin_0/tmux_2to1_3/A
+ tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G
+ tmux_7therm_to_3bin_0/R1/R1 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin tmux_7therm_to_3bin_0/buffer_2/inv_1/vin
+ tmux_7therm_to_3bin_0/R1/m1_n100_n100# tmux_7therm_to_3bin_0/buffer_1/out tmux_7therm_to_3bin_0/buffer_8/in
+ vdd vss tmux_7therm_to_3bin_0/buffer_7/in tmux_7therm_to_3bin_0/buffer_4/out tmux_7therm_to_3bin
C0 comp_p_2/tail vdd 0.00168f
C1 vin comp_p_3/tail 0.00233f
C2 d5 comp_p_3/out_left 0.02324f
C3 comp_p_3/latch_left comp_p_3/vinn 0.00666f
C4 comp_p_4/latch_left comp_p_6/vinn 0.00606f
C5 d1 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0.00131f
C6 comp_p_5/latch_left d6 0.00183f
C7 comp_p_2/latch_left comp_p_0/out_left 0.01472f
C8 vref comp_p_6/vinn 0.00148f
C9 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d3 0
C10 d5 tmux_7therm_to_3bin_0/buffer_5/out 0
C11 comp_p_1/vinn comp_p_0/latch_right 0.1958f
C12 d4 tmux_7therm_to_3bin_0/buffer_0/out 0
C13 vdd d2 1.1602f
C14 vin comp_p_4/tail 0.01181f
C15 tmux_7therm_to_3bin_0/buffer_1/out d2 0
C16 comp_p_4/latch_right d4 0
C17 vbias_generation_0/XR_bias_4/R1 comp_p_4/latch_left 0
C18 vdd tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C19 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vdd 0.00104f
C20 vin comp_p_1/out_left 0.07139f
C21 d0 tmux_7therm_to_3bin_0/buffer_0/out 0
C22 comp_p_5/vinn comp_p_4/tail 0.10856f
C23 comp_p_6/out_left vdd 1.84652f
C24 tmux_7therm_to_3bin_0/R1/R1 vdd 0.00399f
C25 tmux_7therm_to_3bin_0/R1/R1 tmux_7therm_to_3bin_0/buffer_1/out 0
C26 d1 comp_p_3/vinn 0
C27 d6 d2 0.05303f
C28 comp_p_1/vinn d2 0.00152f
C29 vdd tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0.00196f
C30 tmux_7therm_to_3bin_0/buffer_2/out d3 0
C31 vin d1 0.63586f
C32 comp_p_4/out_left comp_p_6/vinn 0.04948f
C33 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d6 0
C34 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin d6 0
C35 dout0 dout1 -0
C36 d1 comp_p_1/tail 0.00457f
C37 comp_p_4/latch_right comp_p_4/vinn 0.00144f
C38 d5 tmux_7therm_to_3bin_0/buffer_0/out 0
C39 vbias_generation_0/XR_bias_4/R1 comp_p_4/out_left 0
C40 tmux_7therm_to_3bin_0/tmux_2to1_3/A vdd 0.00153f
C41 d6 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C42 vdd comp_p_5/latch_right 1.9557f
C43 comp_p_0/latch_left vin 0.00334f
C44 vdd comp_p_3/vinn 1.48772f
C45 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d1 0.00482f
C46 vin vdd 10.39915f
C47 vbias_generation_0/bias_n comp_p_6/vinn 0.43753f
C48 comp_p_0/vinn comp_p_2/out_left 0.0271f
C49 d4 d0 0.03391f
C50 d4 comp_p_5/tail 0.00264f
C51 vdd comp_p_1/tail 0.35563f
C52 comp_p_5/vinn vdd 1.45079f
C53 comp_p_5/latch_right d6 0
C54 comp_p_3/latch_right d2 0.09517f
C55 comp_p_2/vinn comp_p_3/out_left 0
C56 comp_p_3/vinn d6 0
C57 comp_p_1/vinn comp_p_3/vinn 0.03321f
C58 vin vbias_generation_0/XR_bias_2/R2 0.50675f
C59 vin d6 0.01178f
C60 d4 comp_p_4/vinn -0
C61 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d2 0.00483f
C62 vin comp_p_1/vinn 0.97735f
C63 d1 tmux_7therm_to_3bin_0/buffer_2/out 0.00551f
C64 d5 d4 4.51321f
C65 comp_p_2/tail comp_p_3/out_left 0
C66 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin vdd 0
C67 d6 comp_p_1/tail 0
C68 comp_p_5/vinn d6 0.00513f
C69 vin comp_p_6/tail 0
C70 comp_p_6/out_left comp_p_6/vinn 0.14972f
C71 comp_p_5/out_left d3 0.02309f
C72 comp_p_0/vinn comp_p_2/latch_left 0
C73 comp_p_6/vbias_p d3 0
C74 d5 d0 0.04762f
C75 vin comp_p_0/out_left 0.0787f
C76 comp_p_6/latch_left comp_p_5/latch_left 0.00925f
C77 comp_p_3/out_left d2 0.67197f
C78 comp_p_6/vbias_p comp_p_5/out_left -0.0642f
C79 vbias_generation_0/bias_n comp_p_6/latch_left 0.01259f
C80 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d6 0
C81 tmux_7therm_to_3bin_0/R1/R2 d3 0
C82 comp_p_0/vinn comp_p_2/vinn 0.02754f
C83 comp_p_0/vinn comp_p_0/latch_right 0.00236f
C84 comp_p_3/latch_left d3 0
C85 comp_p_3/latch_right comp_p_3/vinn 0.00805f
C86 comp_p_4/latch_right comp_p_5/latch_left 0.02598f
C87 comp_p_5/out_left comp_p_4/tail 0
C88 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d4 0.00384f
C89 comp_p_6/vbias_p comp_p_4/tail 0.31443f
C90 vin comp_p_6/vinn 1.01745f
C91 vbias_generation_0/bias_n comp_p_4/latch_right 0
C92 comp_p_2/vinn comp_p_2/latch_right 0
C93 comp_p_1/out_left d3 0
C94 comp_p_2/latch_right comp_p_0/latch_right 0.01494f
C95 comp_p_1/latch_left d3 0
C96 comp_p_1/latch_right d3 0.00104f
C97 comp_p_6/vbias_p comp_p_1/out_left -0.065f
C98 comp_p_4/latch_left comp_p_4/vinn 0.00288f
C99 comp_p_5/vinn comp_p_6/vinn 0.03037f
C100 vdd tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0.00122f
C101 d2 tmux_7therm_to_3bin_0/buffer_0/out 0
C102 vin vbias_generation_0/XR_bias_4/R1 0.00472f
C103 d1 d3 0.11517f
C104 comp_p_3/out_left comp_p_3/vinn 0.20126f
C105 vin comp_p_3/out_left 0.05071f
C106 comp_p_6/vbias_p d1 0.37529f
C107 comp_p_2/latch_right d2 0.00137f
C108 comp_p_5/latch_left d4 0.06545f
C109 vin comp_p_0/tail 0.01181f
C110 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d6 0.00531f
C111 comp_p_1/latch_left comp_p_3/latch_left 0.00925f
C112 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d5 0.00186f
C113 vbias_generation_0/bias_n d4 0.00802f
C114 comp_p_4/vinn comp_p_4/out_left 0.02516f
C115 comp_p_3/latch_left d1 0
C116 vdd comp_p_6/latch_right 1.95582f
C117 vdd d3 2.3721f
C118 comp_p_6/vbias_p comp_p_0/latch_left 0.37827f
C119 vin comp_p_6/latch_left 0.00266f
C120 comp_p_5/out_left vdd 1.8042f
C121 tmux_7therm_to_3bin_0/buffer_1/out d3 0
C122 comp_p_6/vbias_p vdd 12.48384f
C123 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G d0 0
C124 d4 d2 0.04942f
C125 comp_p_1/out_left d1 0.67001f
C126 comp_p_0/vinn comp_p_3/vinn 0.53686f
C127 d1 comp_p_1/latch_right 0.09536f
C128 comp_p_1/latch_left d1 0.09502f
C129 d4 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C130 comp_p_0/vinn vin 0.81463f
C131 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d4 0.00318f
C132 comp_p_2/out_left comp_p_4/out_left 0.01584f
C133 d3 d6 0.07956f
C134 d0 d2 0.03281f
C135 comp_p_1/vinn d3 0
C136 comp_p_5/out_left d6 0
C137 comp_p_3/tail vdd 0.35691f
C138 comp_p_6/vbias_p vbias_generation_0/XR_bias_2/R2 0.02749f
C139 tmux_7therm_to_3bin_0/R1/R1 d4 0
C140 comp_p_6/out_left d4 0.27385f
C141 vin comp_p_4/latch_right 0.21628f
C142 comp_p_3/latch_left vdd 2.04611f
C143 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vdd 0
C144 comp_p_6/vbias_p comp_p_1/vinn 0.38594f
C145 comp_p_2/latch_right comp_p_3/vinn 0.17593f
C146 vin comp_p_2/latch_right 0.21614f
C147 vdd comp_p_4/tail 0.00166f
C148 d4 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C149 tmux_7therm_to_3bin_0/R1/R1 d0 0.00538f
C150 comp_p_4/latch_right comp_p_5/vinn 0.20935f
C151 comp_p_1/out_left vdd 1.79183f
C152 vdd tmux_7therm_to_3bin_0/buffer_4/out 0.00846f
C153 comp_p_2/out_left comp_p_2/vinn 0.0232f
C154 comp_p_3/tail d6 0
C155 comp_p_6/vbias_p comp_p_0/out_left 0.68459f
C156 d0 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0.00746f
C157 comp_p_1/latch_left vdd 2.04615f
C158 comp_p_1/latch_right vdd 1.96641f
C159 comp_p_3/latch_left d6 0
C160 d5 d2 0.04508f
C161 vbias_generation_0/bias_n comp_p_4/latch_left 0
C162 d1 vdd 1.15842f
C163 d4 comp_p_5/latch_right 0.06539f
C164 d5 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C165 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d5 0
C166 d1 tmux_7therm_to_3bin_0/buffer_1/out 0.01311f
C167 d4 comp_p_3/vinn 0
C168 comp_p_1/out_left d6 0
C169 tmux_7therm_to_3bin_0/tmux_2to1_3/A d0 0
C170 comp_p_1/out_left comp_p_1/vinn 0.19389f
C171 tmux_7therm_to_3bin_0/buffer_4/out d6 0
C172 vin d4 0.72855f
C173 comp_p_1/latch_right d6 0.00271f
C174 comp_p_1/latch_left d6 0
C175 comp_p_1/latch_left comp_p_1/vinn 0.0067f
C176 comp_p_1/latch_right comp_p_1/vinn 0.00799f
C177 comp_p_3/latch_right d3 0.0057f
C178 d5 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C179 comp_p_6/latch_right comp_p_6/vinn 0.00296f
C180 d4 comp_p_1/tail 0
C181 vbias_generation_0/XR_bias_3/R2 comp_p_6/out_left 0.00563f
C182 comp_p_5/vinn d4 0.25734f
C183 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d3 0
C184 d1 d6 0.09f
C185 d1 comp_p_1/vinn 0.26331f
C186 comp_p_6/vbias_p comp_p_6/vinn 0.31983f
C187 comp_p_0/latch_left vdd 0
C188 comp_p_2/vinn comp_p_2/latch_left 0
C189 vin comp_p_5/tail 0.00233f
C190 comp_p_6/vbias_p vbias_generation_0/XR_bias_4/R1 0.02724f
C191 comp_p_3/vinn comp_p_4/vinn 0
C192 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d4 0
C193 comp_p_5/out_left comp_p_3/out_left 0.01584f
C194 vin comp_p_4/vinn 0.52728f
C195 comp_p_6/vbias_p comp_p_3/out_left -0.06014f
C196 d5 comp_p_3/vinn 0
C197 comp_p_0/latch_left comp_p_1/vinn 0.15776f
C198 d5 vin 0.0056f
C199 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d0 0
C200 vdd d6 5.14819f
C201 tmux_7therm_to_3bin_0/R1/m1_n100_n100# d3 0
C202 comp_p_5/vinn comp_p_4/vinn 0.32186f
C203 vdd comp_p_1/vinn 1.45687f
C204 comp_p_6/vbias_p comp_p_0/tail 0.31443f
C205 vbias_generation_0/XR_bias_3/R2 vin 0.08368f
C206 d5 comp_p_1/tail 0
C207 comp_p_3/latch_right comp_p_1/latch_right 0.00925f
C208 comp_p_6/tail vdd 0.35623f
C209 comp_p_2/tail comp_p_2/vinn 0
C210 comp_p_2/out_left comp_p_3/vinn 0.01462f
C211 d4 tmux_7therm_to_3bin_0/buffer_2/out 0
C212 comp_p_2/out_left vin 0.0842f
C213 vin comp_p_4/latch_left 0.00664f
C214 comp_p_3/latch_right d1 0
C215 vdd comp_p_0/out_left 0.01217f
C216 comp_p_0/latch_right d2 0.01472f
C217 comp_p_1/vinn d6 0
C218 vin vref 0.03789f
C219 d1 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0.00173f
C220 d5 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C221 comp_p_5/vinn comp_p_4/latch_left 0.16266f
C222 d3 tmux_7therm_to_3bin_0/buffer_0/out 0
C223 comp_p_2/tail d2 -0.00224f
C224 comp_p_0/vinn comp_p_6/vbias_p 0.12305f
C225 comp_p_0/tail comp_p_1/out_left 0
C226 comp_p_1/vinn comp_p_0/out_left 0.04644f
C227 vbias_generation_0/bias_n comp_p_6/out_left 0.00925f
C228 comp_p_5/out_left comp_p_4/latch_right 0
C229 d4 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0.00248f
C230 comp_p_6/vbias_p comp_p_4/latch_right 0.40389f
C231 comp_p_3/latch_right vdd 1.95698f
C232 vdd tmux_7therm_to_3bin_0/buffer_7/in 0.0027f
C233 comp_p_2/latch_left comp_p_3/vinn 0.15548f
C234 vin comp_p_4/out_left 0.0859f
C235 comp_p_6/vbias_p comp_p_2/latch_right 0.40389f
C236 vdd comp_p_6/vinn 1.11418f
C237 vin comp_p_2/latch_left 0.00664f
C238 comp_p_0/tail d1 -0.00224f
C239 comp_p_5/vinn comp_p_4/out_left 0.01843f
C240 tmux_7therm_to_3bin_0/R1/R1 d2 0.00763f
C241 tmux_7therm_to_3bin_0/buffer_6/out d6 0
C242 comp_p_3/latch_right d6 0.00265f
C243 d2 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C244 comp_p_2/vinn comp_p_3/vinn 0.31389f
C245 comp_p_0/vinn comp_p_1/out_left 0
C246 vbias_generation_0/XR_bias_2/R2 comp_p_6/vinn 0.00358f
C247 comp_p_3/out_left vdd 1.79594f
C248 comp_p_3/latch_left comp_p_2/latch_right 0.02598f
C249 vin comp_p_2/vinn 0.52215f
C250 vin comp_p_0/latch_right 0.21598f
C251 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d6 0
C252 d4 comp_p_6/latch_right 0.06065f
C253 d4 d3 2.88908f
C254 vbias_generation_0/bias_n vin 0.0214f
C255 comp_p_5/out_left d4 0.61081f
C256 d5 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0
C257 comp_p_6/vbias_p d4 0.37293f
C258 comp_p_5/latch_left comp_p_5/vinn 0.00674f
C259 comp_p_0/tail vdd 0.00166f
C260 comp_p_2/tail comp_p_3/vinn 0.14685f
C261 comp_p_0/vinn d1 -0
C262 comp_p_2/tail vin 0.0104f
C263 d0 d3 0.03225f
C264 d1 tmux_7therm_to_3bin_0/buffer_0/out 0
C265 comp_p_6/vbias_p d0 0.00465f
C266 comp_p_3/out_left d6 0
C267 comp_p_3/vinn d2 0.24742f
C268 vin d2 0.72189f
C269 comp_p_6/latch_left vdd 2.04625f
C270 comp_p_3/tail d4 0
C271 d1 comp_p_2/latch_right 0.01472f
C272 comp_p_3/latch_left d4 0
C273 comp_p_0/tail comp_p_1/vinn 0.10698f
C274 comp_p_1/tail d2 0
C275 d4 comp_p_4/tail -0.00224f
C276 comp_p_0/vinn comp_p_0/latch_left 0.02494f
C277 comp_p_5/out_left comp_p_4/vinn 0
C278 vin comp_p_6/out_left 0.06197f
C279 comp_p_6/vbias_p comp_p_4/vinn 0.12306f
C280 d5 d3 0.16529f
C281 comp_p_0/vinn vdd 0.01961f
C282 comp_p_1/out_left d4 0
C283 d5 comp_p_5/out_left 0
C284 vdd tmux_7therm_to_3bin_0/buffer_0/out 0
C285 comp_p_6/vbias_p d5 0
C286 d4 tmux_7therm_to_3bin_0/buffer_4/out 0
C287 comp_p_1/latch_right d4 0
C288 comp_p_1/latch_left d4 0
C289 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vdd 0.00166f
C290 comp_p_4/latch_right vdd 0.00589f
C291 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d2 0.00171f
C292 comp_p_1/out_left d0 -0
C293 comp_p_2/latch_right vdd 0.00592f
C294 d1 d4 0.33457f
C295 comp_p_0/vinn comp_p_1/vinn 0.94729f
C296 d5 comp_p_3/tail 0
C297 comp_p_6/vbias_p comp_p_2/out_left 0.68901f
C298 d6 tmux_7therm_to_3bin_0/buffer_0/out 0
C299 vbias_generation_0/XR_bias_4/R1 comp_p_6/vinn 0.51064f
C300 comp_p_6/vbias_p comp_p_4/latch_left 0.37827f
C301 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin tmux_7therm_to_3bin_0/R1/R1 0
C302 d5 comp_p_3/latch_left 0
C303 d1 d0 1.12322f
C304 vin comp_p_3/vinn 0.65736f
C305 comp_p_2/latch_right comp_p_1/vinn 0.00771f
C306 tmux_7therm_to_3bin_0/buffer_2/out d2 0
C307 comp_p_5/vinn comp_p_5/latch_right 0.00802f
C308 comp_p_0/vinn comp_p_0/out_left 0.02276f
C309 d5 comp_p_1/out_left 0
C310 comp_p_5/vinn comp_p_3/vinn 0.0226f
C311 d5 tmux_7therm_to_3bin_0/buffer_4/out 0
C312 d5 comp_p_1/latch_right 0.0019f
C313 d5 comp_p_1/latch_left 0
C314 vin comp_p_1/tail 0.00233f
C315 d4 vdd 1.46527f
C316 vin comp_p_5/vinn 0.66275f
C317 d4 tmux_7therm_to_3bin_0/buffer_1/out 0
C318 d5 d1 0.26099f
C319 vdd d0 2.71992f
C320 comp_p_6/latch_left comp_p_6/vinn 0.00473f
C321 comp_p_6/vbias_p comp_p_4/out_left 0.69034f
C322 comp_p_6/vbias_p comp_p_2/latch_left 0.37827f
C323 vdd comp_p_5/tail 0.35567f
C324 d4 d6 0.79887f
C325 d4 comp_p_1/vinn 0
C326 comp_p_6/tail d4 0.00252f
C327 d0 d6 0.09283f
C328 vdd comp_p_4/vinn 0.03662f
C329 vbias_generation_0/bias_n comp_p_6/latch_right 0
C330 comp_p_6/vbias_p comp_p_2/vinn 0.12413f
C331 comp_p_4/latch_right comp_p_6/vinn 0.00583f
C332 comp_p_6/vbias_p comp_p_0/latch_right 0.40389f
C333 d5 vdd 2.33637f
C334 d6 comp_p_5/tail 0
C335 comp_p_6/vbias_p vbias_generation_0/bias_n 0
C336 vbias_generation_0/XR_bias_3/R2 vdd 0.08059f
C337 comp_p_6/vbias_p comp_p_2/tail 0.31443f
C338 comp_p_4/latch_right vbias_generation_0/XR_bias_4/R1 0
C339 comp_p_0/latch_left comp_p_2/out_left 0.01472f
C340 d3 d2 2.50136f
C341 comp_p_2/out_left vdd 0.02487f
C342 vdd comp_p_4/latch_left 0
C343 d5 d6 4.44886f
C344 comp_p_6/vbias_p d2 0.37534f
C345 d5 comp_p_1/vinn 0
C346 tmux_7therm_to_3bin_0/buffer_6/out d4 0.013f
C347 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d3 0
C348 comp_p_3/out_left comp_p_2/latch_right 0
C349 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin d3 0.00238f
C350 vdd vref 0
C351 comp_p_3/latch_right d4 0.00133f
C352 tmux_7therm_to_3bin_0/R1/R1 d3 0
C353 comp_p_1/out_left comp_p_0/latch_right 0
C354 d4 comp_p_6/vinn 0.06841f
C355 comp_p_6/vbias_p comp_p_6/out_left -0.05282f
C356 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d4 0
C357 comp_p_1/latch_left comp_p_0/latch_right 0.02598f
C358 d3 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C359 vbias_generation_0/XR_bias_3/R2 comp_p_6/tail 0
C360 comp_p_3/tail d2 0.00272f
C361 comp_p_2/out_left comp_p_1/vinn 0.00265f
C362 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin vdd 0.00104f
C363 comp_p_3/latch_left d2 0.09614f
C364 d1 comp_p_0/latch_right 0
C365 comp_p_0/latch_left comp_p_2/latch_left 0.01494f
C366 vdd comp_p_4/out_left 0.02489f
C367 comp_p_3/out_left d4 0
C368 comp_p_2/latch_left vdd 0
C369 comp_p_1/out_left d2 0
C370 comp_p_2/out_left comp_p_0/out_left 0.09264f
C371 comp_p_5/latch_right comp_p_6/latch_right 0.00925f
C372 tmux_7therm_to_3bin_0/buffer_5/out d4 0.01353f
C373 comp_p_1/latch_right d2 0.00123f
C374 comp_p_1/latch_left d2 0
C375 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d6 0
C376 comp_p_3/vinn d3 0.0076f
C377 d5 comp_p_3/latch_right 0.00185f
C378 vin d3 0.00158f
C379 comp_p_6/vbias_p comp_p_3/vinn 0.38072f
C380 vin comp_p_5/out_left 0.06043f
C381 d1 d2 3.44306f
C382 comp_p_5/latch_left vdd 2.0461f
C383 comp_p_6/vbias_p vin 1.44761f
C384 d5 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C385 comp_p_2/vinn vdd 0.04727f
C386 vdd comp_p_0/latch_right 0.00588f
C387 comp_p_2/latch_left comp_p_1/vinn 0.01672f
C388 d3 comp_p_1/tail 0
C389 vbias_generation_0/bias_n vdd 0.0189f
C390 comp_p_6/latch_left d4 0.06068f
C391 vbias_generation_0/XR_bias_3/R2 comp_p_6/vinn 0.06411f
C392 comp_p_5/out_left comp_p_5/vinn 0.19629f
C393 tmux_7therm_to_3bin_0/buffer_8/in vdd 0
C394 comp_p_6/vbias_p comp_p_5/vinn 0.407f
C395 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G vdd 0.00166f
C396 d1 tmux_7therm_to_3bin_0/R1/R1 0.00785f
C397 tmux_7therm_to_3bin_0/tmux_2to1_3/A vss 0.4939f
C398 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G vss 0.55051f
C399 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin vss 0.52606f
C400 dout2 vss 0.32356f
C401 tmux_7therm_to_3bin_0/buffer_8/inv_1/vin vss 0.52606f
C402 dout1 vss 0.32356f
C403 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vss 0.52606f
C404 dout0 vss 0.32356f
C405 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin vss 0.52765f
C406 tmux_7therm_to_3bin_0/buffer_6/out vss 0.67609f
C407 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin vss 0.52606f
C408 tmux_7therm_to_3bin_0/buffer_5/out vss 0.70857f
C409 vdd vss 0.3833p
C410 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vss 0.52606f
C411 tmux_7therm_to_3bin_0/buffer_4/out vss 0.70167f
C412 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin vss 0.52606f
C413 tmux_7therm_to_3bin_0/R1/R2 vss 0.22083f
C414 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin vss 0.52811f
C415 tmux_7therm_to_3bin_0/buffer_2/out vss 0.28552f
C416 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin vss 0.52606f
C417 tmux_7therm_to_3bin_0/buffer_1/out vss 0.30295f
C418 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin vss 0.52606f
C419 tmux_7therm_to_3bin_0/buffer_0/out vss 0.30577f
C420 tmux_7therm_to_3bin_0/R1/m1_n100_n100# vss 0.10692f
C421 tmux_7therm_to_3bin_0/buffer_8/in vss 1.28735f
C422 tmux_7therm_to_3bin_0/buffer_7/in vss 0.74661f
C423 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vss 0.55051f
C424 tmux_7therm_to_3bin_0/R1/R1 vss 3.00001f
C425 tmux_7therm_to_3bin_0/tmux_2to1_3/B vss 0.41874f
C426 tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G vss 0.55051f
C427 tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G vss 0.55051f
C428 vin vss 20.78606f
C429 comp_p_6/tail vss 1.09633f
C430 d6 vss 4.91925f
C431 comp_p_6/latch_right vss 3.49411f
C432 comp_p_6/out_left vss 2.08947f
C433 comp_p_6/latch_left vss 3.68918f
C434 comp_p_5/tail vss 1.09613f
C435 d5 vss 3.00569f
C436 comp_p_5/latch_right vss 3.49805f
C437 comp_p_5/out_left vss 2.08667f
C438 comp_p_5/latch_left vss 3.68855f
C439 comp_p_4/tail vss 1.56897f
C440 d4 vss 9.4397f
C441 comp_p_4/latch_right vss 5.50989f
C442 comp_p_4/out_left vss 4.34925f
C443 comp_p_4/latch_left vss 6.03696f
C444 comp_p_3/tail vss 1.09611f
C445 d3 vss 2.71104f
C446 comp_p_3/latch_right vss 3.5009f
C447 comp_p_3/out_left vss 2.06137f
C448 comp_p_3/latch_left vss 3.68751f
C449 comp_p_2/tail vss 1.56898f
C450 d2 vss 7.1799f
C451 comp_p_2/latch_right vss 5.49653f
C452 comp_p_2/out_left vss 4.34035f
C453 comp_p_2/latch_left vss 6.03407f
C454 comp_p_0/tail vss 1.56897f
C455 d1 vss 7.38418f
C456 comp_p_0/latch_right vss 5.50255f
C457 comp_p_0/out_left vss 4.40824f
C458 comp_p_0/latch_left vss 6.03535f
C459 comp_p_1/tail vss 1.09611f
C460 d0 vss 2.80029f
C461 comp_p_1/latch_right vss 3.49227f
C462 comp_p_1/out_left vss 2.0627f
C463 comp_p_1/latch_left vss 3.68751f
C464 comp_p_0/vinn vss 6.06348f
C465 comp_p_2/vinn vss 4.46291f
C466 comp_p_3/vinn vss 7.47636f
C467 comp_p_4/vinn vss 4.49649f
C468 comp_p_5/vinn vss 7.17599f
C469 comp_p_6/vinn vss 8.16656f
C470 comp_p_1/vinn vss 8.18212f
C471 vref vss 4.52985f
C472 vbias_generation_0/bias_n vss 2.63421f
C473 vbias_generation_0/XR_bias_4/R1 vss 1.61917f
C474 vbias_generation_0/XR_bias_3/R2 vss 1.9113f
C475 vbias_generation_0/XR_bias_2/R2 vss 1.5274f
C476 comp_p_6/vbias_p vss 14.49086f
.ends

.subckt tt_um_tinyflash_extracted clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND
XflashADC_3bit_0 uo_out[0] uo_out[1] uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out
+ flashADC_3bit_0/vbias_generation_0/bias_n flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin flashADC_3bit_0/comp_p_3/latch_left
+ flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in
+ flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in
+ flashADC_3bit_0/comp_p_5/latch_left flashADC_3bit_0/vbias_generation_0/XR_bias_2/R2
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/m1_n100_n100# flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin
+ flashADC_3bit_0/comp_p_6/latch_left flashADC_3bit_0/comp_p_1/out_left flashADC_3bit_0/comp_p_6/tail
+ flashADC_3bit_0/comp_p_0/latch_right flashADC_3bit_0/comp_p_1/latch_right flashADC_3bit_0/comp_p_2/latch_right
+ flashADC_3bit_0/comp_p_3/latch_right flashADC_3bit_0/comp_p_3/tail flashADC_3bit_0/comp_p_4/latch_right
+ flashADC_3bit_0/comp_p_5/latch_right flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out flashADC_3bit_0/comp_p_4/out_left
+ flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_6/latch_right flashADC_3bit_0/comp_p_0/tail
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 flashADC_3bit_0/comp_p_2/latch_left
+ flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G
+ uo_out[4] flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G
+ flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out
+ flashADC_3bit_0/comp_p_0/out_left flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G flashADC_3bit_0/comp_p_6/vinn
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out uo_out[5] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin
+ flashADC_3bit_0/comp_p_4/tail flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/comp_p_0/latch_left
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin
+ uo_out[7] flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B
+ flashADC_3bit_0/comp_p_1/tail flashADC_3bit_0/comp_p_0/vinn ua[0] flashADC_3bit_0/comp_p_6/out_left
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A flashADC_3bit_0/comp_p_1/latch_left
+ VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out uio_out[0] uo_out[6] uo_out[3]
+ flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_2/vinn ua[1] flashADC_3bit_0/comp_p_5/out_left
+ flashADC_3bit_0/vbias_generation_0/XR_bias_3/R2 uio_out[1] VGND flashADC_3bit_0/comp_p_3/out_left
+ flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit
X0 flashADC_3bit_0/comp_p_0/tail ua[0].t7 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X1 flashADC_3bit_0/comp_p_6/tail ua[0].t25 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X2 flashADC_3bit_0/comp_p_0/latch_left flashADC_3bit_0/comp_p_0/latch_right.t2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X3 uo_out[4] flashADC_3bit_0/comp_p_0/latch_right.t3 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X4 flashADC_3bit_0/comp_p_4/tail ua[0].t16 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X5 flashADC_3bit_0/comp_p_2/tail ua[0].t9 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X6 flashADC_3bit_0/comp_p_5/tail ua[0].t22 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X7 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin uo_out[6].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X8 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin uo_out[5].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X9 flashADC_3bit_0/comp_p_2/tail ua[0].t8 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X10 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin uio_out[0].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X11 flashADC_3bit_0/comp_p_1/tail ua[0].t0 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X12 flashADC_3bit_0/comp_p_3/tail ua[0].t15 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X13 flashADC_3bit_0/comp_p_4/tail ua[0].t17 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X14 flashADC_3bit_0/comp_p_5/tail ua[0].t23 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X15 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin uio_out[1].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X16 flashADC_3bit_0/comp_p_1/tail ua[0].t1 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X17 flashADC_3bit_0/comp_p_6/tail ua[0].t27 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X18 flashADC_3bit_0/comp_p_6/out_left flashADC_3bit_0/comp_p_6/latch_left.t3 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X19 flashADC_3bit_0/comp_p_6/tail ua[0].t26 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X20 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin uo_out[4].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X21 VDPWR flashADC_3bit_0/comp_p_0/out_left.t0 flashADC_3bit_0/comp_p_0/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X22 flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/comp_p_2/latch_left.t3 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X23 VDPWR flashADC_3bit_0/comp_p_5/out_left.t0 flashADC_3bit_0/comp_p_5/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X24 flashADC_3bit_0/comp_p_4/tail ua[0].t18 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X25 VDPWR flashADC_3bit_0/comp_p_5/out_left.t2 uio_out[0] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X26 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X27 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin uo_out[7].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X28 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin uio_out[1].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X29 flashADC_3bit_0/comp_p_0/tail ua[0].t4 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X30 flashADC_3bit_0/comp_p_1/tail ua[0].t2 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X31 flashADC_3bit_0/comp_p_2/tail ua[0].t11 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X32 flashADC_3bit_0/comp_p_3/tail ua[0].t14 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X33 flashADC_3bit_0/comp_p_4/latch_left.t1 flashADC_3bit_0/comp_p_4/latch_left.t0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X34 flashADC_3bit_0/comp_p_4/tail ua[0].t19 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X35 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin uo_out[6].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X36 flashADC_3bit_0/comp_p_0/tail ua[0].t5 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X37 flashADC_3bit_0/comp_p_1/tail ua[0].t3 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X38 flashADC_3bit_0/comp_p_4/out_left flashADC_3bit_0/comp_p_4/latch_left.t3 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X39 flashADC_3bit_0/comp_p_6/tail ua[0].t24 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X40 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin uio_out[0].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X41 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin uo_out[5].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X42 flashADC_3bit_0/comp_p_0/latch_right.t1 flashADC_3bit_0/comp_p_0/latch_right.t0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X43 flashADC_3bit_0/comp_p_5/tail ua[0].t20 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X44 flashADC_3bit_0/comp_p_2/latch_left.t1 flashADC_3bit_0/comp_p_2/latch_left.t0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X45 flashADC_3bit_0/comp_p_3/tail ua[0].t13 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X46 flashADC_3bit_0/comp_p_4/latch_right flashADC_3bit_0/comp_p_4/latch_left.t2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X47 flashADC_3bit_0/comp_p_6/latch_left.t1 flashADC_3bit_0/comp_p_6/latch_left.t0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X48 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin uo_out[7].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X49 VDPWR flashADC_3bit_0/comp_p_1/out_left.t0 flashADC_3bit_0/comp_p_1/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X50 flashADC_3bit_0/comp_p_3/tail ua[0].t12 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X51 VDPWR flashADC_3bit_0/comp_p_1/out_left.t2 uo_out[3] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X52 VDPWR flashADC_3bit_0/comp_p_0/out_left.t2 uo_out[4] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X53 flashADC_3bit_0/comp_p_5/tail ua[0].t21 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X54 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin uo_out[4].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X55 flashADC_3bit_0/comp_p_0/tail ua[0].t6 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X56 flashADC_3bit_0/comp_p_2/tail ua[0].t10 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X57 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X58 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_2/latch_left.t2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X59 flashADC_3bit_0/comp_p_6/latch_right flashADC_3bit_0/comp_p_6/latch_left.t2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
R0 VGND.n952 VGND.n951 28249.5
R1 VGND.n606 VGND.n16 15045.2
R2 VGND.n351 VGND.n15 12367.9
R3 VGND.n15 VGND.n14 12039.7
R4 VGND.n953 VGND.n952 11644.9
R5 VGND.n607 VGND.n606 11496.8
R6 VGND.n968 VGND.n965 10655.8
R7 VGND.n354 VGND.n349 10261.4
R8 VGND.n352 VGND.n349 10261.4
R9 VGND.n950 VGND.n267 10261.4
R10 VGND.n950 VGND.n268 10261.4
R11 VGND.n156 VGND.n153 8494.18
R12 VGND.n175 VGND.n137 8494.18
R13 VGND.n175 VGND.n174 8494.18
R14 VGND.n1023 VGND.n1022 7442.95
R15 VGND.n161 VGND.n160 7120.97
R16 VGND.n160 VGND.n148 7120.97
R17 VGND.n166 VGND.n142 7120.97
R18 VGND.n166 VGND.n165 7120.97
R19 VGND.n172 VGND.n139 7120.97
R20 VGND.n173 VGND.n172 7120.97
R21 VGND.n608 VGND.n265 6402.87
R22 VGND.n364 VGND.n344 6385.12
R23 VGND.n344 VGND.n342 6385.12
R24 VGND.n359 VGND.n345 6385.12
R25 VGND.n359 VGND.n358 6385.12
R26 VGND.n369 VGND.n336 6385.12
R27 VGND.n369 VGND.n368 6385.12
R28 VGND.n376 VGND.n333 6385.12
R29 VGND.n377 VGND.n376 6385.12
R30 VGND.n385 VGND.n321 6385.12
R31 VGND.n321 VGND.n319 6385.12
R32 VGND.n381 VGND.n322 6385.12
R33 VGND.n381 VGND.n326 6385.12
R34 VGND.n390 VGND.n300 6385.12
R35 VGND.n390 VGND.n389 6385.12
R36 VGND.n306 VGND.n299 6385.12
R37 VGND.n307 VGND.n306 6385.12
R38 VGND.n310 VGND.n309 6385.12
R39 VGND.n310 VGND.n305 6385.12
R40 VGND.n1026 VGND.n8 5440.68
R41 VGND.n45 VGND.n35 5440.68
R42 VGND.n1004 VGND.n33 5440.68
R43 VGND.n292 VGND.n282 5440.68
R44 VGND.n645 VGND.n451 5440.68
R45 VGND.n427 VGND.n283 5440.68
R46 VGND.n655 VGND.n452 5440.68
R47 VGND.n233 VGND.n182 5255.26
R48 VGND.n81 VGND.n69 5255.26
R49 VGND.n91 VGND.n70 5255.26
R50 VGND.n435 VGND.n408 5255.26
R51 VGND.n637 VGND.n474 5255.26
R52 VGND.n716 VGND.n409 5255.26
R53 VGND.n616 VGND.n475 5255.26
R54 VGND.n236 VGND.n179 5116.21
R55 VGND.n236 VGND.n135 5116.21
R56 VGND.n240 VGND.n179 5116.21
R57 VGND.n240 VGND.n135 5116.21
R58 VGND.n207 VGND.n185 4536.79
R59 VGND.n219 VGND.n197 4536.79
R60 VGND.n220 VGND.n219 4536.79
R61 VGND.n228 VGND.n185 4536.79
R62 VGND.n119 VGND.n77 4536.79
R63 VGND.n85 VGND.n77 4536.79
R64 VGND.n994 VGND.n46 4536.79
R65 VGND.n996 VGND.n46 4536.79
R66 VGND.n55 VGND.n52 4536.79
R67 VGND.n993 VGND.n55 4536.79
R68 VGND.n87 VGND.n86 4536.79
R69 VGND.n117 VGND.n87 4536.79
R70 VGND.n726 VGND.n415 4536.79
R71 VGND.n417 VGND.n415 4536.79
R72 VGND.n740 VGND.n294 4536.79
R73 VGND.n742 VGND.n294 4536.79
R74 VGND.n667 VGND.n481 4536.79
R75 VGND.n610 VGND.n481 4536.79
R76 VGND.n682 VGND.n462 4536.79
R77 VGND.n463 VGND.n462 4536.79
R78 VGND.n399 VGND.n295 4536.79
R79 VGND.n739 VGND.n399 4536.79
R80 VGND.n419 VGND.n418 4536.79
R81 VGND.n724 VGND.n419 4536.79
R82 VGND.n467 VGND.n464 4536.79
R83 VGND.n680 VGND.n467 4536.79
R84 VGND.n612 VGND.n611 4536.79
R85 VGND.n665 VGND.n612 4536.79
R86 VGND.n1021 VGND.n16 4301.43
R87 VGND.n233 VGND.n7 4131.21
R88 VGND.n210 VGND.n209 4131.21
R89 VGND.n213 VGND.n212 4131.21
R90 VGND.n226 VGND.n188 4131.21
R91 VGND.n222 VGND.n195 4131.21
R92 VGND.n69 VGND.n68 4131.21
R93 VGND.n123 VGND.n40 4131.21
R94 VGND.n1002 VGND.n41 4131.21
R95 VGND.n125 VGND.n65 4131.21
R96 VGND.n997 VGND.n39 4131.21
R97 VGND.n70 VGND.n32 4131.21
R98 VGND.n104 VGND.n72 4131.21
R99 VGND.n54 VGND.n38 4131.21
R100 VGND.n103 VGND.n71 4131.21
R101 VGND.n107 VGND.n36 4131.21
R102 VGND.n704 VGND.n408 4131.21
R103 VGND.n730 VGND.n287 4131.21
R104 VGND.n748 VGND.n288 4131.21
R105 VGND.n703 VGND.n411 4131.21
R106 VGND.n743 VGND.n286 4131.21
R107 VGND.n640 VGND.n474 4131.21
R108 VGND.n671 VGND.n456 4131.21
R109 VGND.n688 VGND.n457 4131.21
R110 VGND.n477 VGND.n448 4131.21
R111 VGND.n690 VGND.n449 4131.21
R112 VGND.n423 VGND.n409 4131.21
R113 VGND.n732 VGND.n406 4131.21
R114 VGND.n398 VGND.n285 4131.21
R115 VGND.n410 VGND.n279 4131.21
R116 VGND.n750 VGND.n280 4131.21
R117 VGND.n621 VGND.n475 4131.21
R118 VGND.n673 VGND.n472 4131.21
R119 VGND.n466 VGND.n455 4131.21
R120 VGND.n623 VGND.n476 4131.21
R121 VGND.n654 VGND.n453 4131.21
R122 VGND.n543 VGND.n542 4116.13
R123 VGND.n1026 VGND.n7 3945.79
R124 VGND.n209 VGND.n200 3945.79
R125 VGND.n212 VGND.n210 3945.79
R126 VGND.n226 VGND.n186 3945.79
R127 VGND.n222 VGND.n188 3945.79
R128 VGND.n68 VGND.n35 3945.79
R129 VGND.n123 VGND.n73 3945.79
R130 VGND.n1002 VGND.n40 3945.79
R131 VGND.n125 VGND.n63 3945.79
R132 VGND.n65 VGND.n39 3945.79
R133 VGND.n1004 VGND.n32 3945.79
R134 VGND.n93 VGND.n72 3945.79
R135 VGND.n104 VGND.n38 3945.79
R136 VGND.n88 VGND.n71 3945.79
R137 VGND.n103 VGND.n36 3945.79
R138 VGND.n704 VGND.n282 3945.79
R139 VGND.n730 VGND.n412 3945.79
R140 VGND.n748 VGND.n287 3945.79
R141 VGND.n434 VGND.n411 3945.79
R142 VGND.n703 VGND.n286 3945.79
R143 VGND.n640 VGND.n451 3945.79
R144 VGND.n671 VGND.n478 3945.79
R145 VGND.n688 VGND.n456 3945.79
R146 VGND.n636 VGND.n477 3945.79
R147 VGND.n690 VGND.n448 3945.79
R148 VGND.n423 VGND.n283 3945.79
R149 VGND.n732 VGND.n404 3945.79
R150 VGND.n406 VGND.n285 3945.79
R151 VGND.n420 VGND.n410 3945.79
R152 VGND.n750 VGND.n279 3945.79
R153 VGND.n621 VGND.n452 3945.79
R154 VGND.n673 VGND.n471 3945.79
R155 VGND.n472 VGND.n455 3945.79
R156 VGND.n613 VGND.n476 3945.79
R157 VGND.n623 VGND.n453 3945.79
R158 VGND.n389 VGND.n388 3876.26
R159 VGND.n388 VGND.n319 3876.26
R160 VGND.n368 VGND.n367 3876.26
R161 VGND.n367 VGND.n342 3876.26
R162 VGND.n358 VGND.n354 3876.26
R163 VGND.n364 VGND.n363 3876.26
R164 VGND.n363 VGND.n345 3876.26
R165 VGND.n352 VGND.n345 3876.26
R166 VGND.n357 VGND.n342 3876.26
R167 VGND.n358 VGND.n357 3876.26
R168 VGND.n373 VGND.n333 3876.26
R169 VGND.n373 VGND.n336 3876.26
R170 VGND.n365 VGND.n336 3876.26
R171 VGND.n365 VGND.n364 3876.26
R172 VGND.n378 VGND.n326 3876.26
R173 VGND.n378 VGND.n377 3876.26
R174 VGND.n377 VGND.n332 3876.26
R175 VGND.n368 VGND.n332 3876.26
R176 VGND.n385 VGND.n384 3876.26
R177 VGND.n384 VGND.n322 3876.26
R178 VGND.n337 VGND.n322 3876.26
R179 VGND.n337 VGND.n333 3876.26
R180 VGND.n324 VGND.n319 3876.26
R181 VGND.n326 VGND.n324 3876.26
R182 VGND.n394 VGND.n299 3876.26
R183 VGND.n394 VGND.n300 3876.26
R184 VGND.n386 VGND.n300 3876.26
R185 VGND.n386 VGND.n385 3876.26
R186 VGND.n316 VGND.n305 3876.26
R187 VGND.n316 VGND.n307 3876.26
R188 VGND.n307 VGND.n297 3876.26
R189 VGND.n389 VGND.n297 3876.26
R190 VGND.n309 VGND.n267 3876.26
R191 VGND.n314 VGND.n309 3876.26
R192 VGND.n314 VGND.n299 3876.26
R193 VGND.n305 VGND.n268 3876.26
R194 VGND.n952 VGND.n265 3303.94
R195 VGND.n207 VGND.n200 3227.32
R196 VGND.n213 VGND.n197 3227.32
R197 VGND.n228 VGND.n186 3227.32
R198 VGND.n220 VGND.n195 3227.32
R199 VGND.n119 VGND.n73 3227.32
R200 VGND.n994 VGND.n41 3227.32
R201 VGND.n85 VGND.n63 3227.32
R202 VGND.n997 VGND.n996 3227.32
R203 VGND.n93 VGND.n86 3227.32
R204 VGND.n993 VGND.n54 3227.32
R205 VGND.n117 VGND.n88 3227.32
R206 VGND.n107 VGND.n52 3227.32
R207 VGND.n726 VGND.n412 3227.32
R208 VGND.n740 VGND.n288 3227.32
R209 VGND.n434 VGND.n417 3227.32
R210 VGND.n743 VGND.n742 3227.32
R211 VGND.n667 VGND.n478 3227.32
R212 VGND.n682 VGND.n457 3227.32
R213 VGND.n636 VGND.n610 3227.32
R214 VGND.n463 VGND.n449 3227.32
R215 VGND.n418 VGND.n404 3227.32
R216 VGND.n739 VGND.n398 3227.32
R217 VGND.n724 VGND.n420 3227.32
R218 VGND.n295 VGND.n280 3227.32
R219 VGND.n611 VGND.n471 3227.32
R220 VGND.n680 VGND.n466 3227.32
R221 VGND.n665 VGND.n613 3227.32
R222 VGND.n654 VGND.n464 3227.32
R223 VGND.n1022 VGND.n1021 2670.7
R224 VGND.n608 VGND.n607 2649.46
R225 VGND.n591 VGND.n588 2306.06
R226 VGND.n604 VGND.n588 2306.06
R227 VGND.n591 VGND.n589 2306.06
R228 VGND.n604 VGND.n589 2306.06
R229 VGND.n967 VGND.n257 2306.06
R230 VGND.n975 VGND.n257 2306.06
R231 VGND.n967 VGND.n258 2306.06
R232 VGND.n975 VGND.n258 2306.06
R233 VGND.n595 VGND.n594 2306.06
R234 VGND.n594 VGND.n587 2306.06
R235 VGND.n596 VGND.n595 2306.06
R236 VGND.n596 VGND.n587 2306.06
R237 VGND.n963 VGND.n19 2306.06
R238 VGND.n963 VGND.n20 2306.06
R239 VGND.n1019 VGND.n19 2306.06
R240 VGND.n1019 VGND.n20 2306.06
R241 VGND.n961 VGND.n955 2306.06
R242 VGND.n961 VGND.n956 2306.06
R243 VGND.n955 VGND.n18 2306.06
R244 VGND.n956 VGND.n18 2306.06
R245 VGND.n573 VGND.n484 2306.06
R246 VGND.n584 VGND.n484 2306.06
R247 VGND.n573 VGND.n485 2306.06
R248 VGND.n584 VGND.n485 2306.06
R249 VGND.n560 VGND.n491 2306.06
R250 VGND.n570 VGND.n491 2306.06
R251 VGND.n560 VGND.n492 2306.06
R252 VGND.n570 VGND.n492 2306.06
R253 VGND.n547 VGND.n514 2306.06
R254 VGND.n545 VGND.n514 2306.06
R255 VGND.n557 VGND.n499 2306.06
R256 VGND.n557 VGND.n500 2306.06
R257 VGND.n526 VGND.n516 2306.06
R258 VGND.n541 VGND.n516 2306.06
R259 VGND.n526 VGND.n517 2306.06
R260 VGND.n541 VGND.n517 2306.06
R261 VGND.n522 VGND.n520 2306.06
R262 VGND.n529 VGND.n520 2306.06
R263 VGND.n523 VGND.n522 2306.06
R264 VGND.n529 VGND.n523 2306.06
R265 VGND.n575 VGND.n488 2306.06
R266 VGND.n488 VGND.n483 2306.06
R267 VGND.n576 VGND.n575 2306.06
R268 VGND.n576 VGND.n483 2306.06
R269 VGND.n562 VGND.n497 2306.06
R270 VGND.n497 VGND.n490 2306.06
R271 VGND.n563 VGND.n562 2306.06
R272 VGND.n563 VGND.n490 2306.06
R273 VGND.n811 VGND.n793 2306.06
R274 VGND.n802 VGND.n793 2306.06
R275 VGND.n811 VGND.n794 2306.06
R276 VGND.n802 VGND.n794 2306.06
R277 VGND.n821 VGND.n783 2306.06
R278 VGND.n813 VGND.n783 2306.06
R279 VGND.n821 VGND.n784 2306.06
R280 VGND.n813 VGND.n784 2306.06
R281 VGND.n922 VGND.n918 2306.06
R282 VGND.n922 VGND.n919 2306.06
R283 VGND.n932 VGND.n778 2306.06
R284 VGND.n779 VGND.n778 2306.06
R285 VGND.n884 VGND.n858 2306.06
R286 VGND.n899 VGND.n858 2306.06
R287 VGND.n884 VGND.n859 2306.06
R288 VGND.n899 VGND.n859 2306.06
R289 VGND.n868 VGND.n865 2306.06
R290 VGND.n881 VGND.n865 2306.06
R291 VGND.n868 VGND.n866 2306.06
R292 VGND.n881 VGND.n866 2306.06
R293 VGND.n800 VGND.n791 2306.06
R294 VGND.n804 VGND.n800 2306.06
R295 VGND.n801 VGND.n791 2306.06
R296 VGND.n804 VGND.n801 2306.06
R297 VGND.n789 VGND.n781 2306.06
R298 VGND.n815 VGND.n789 2306.06
R299 VGND.n790 VGND.n781 2306.06
R300 VGND.n815 VGND.n790 2306.06
R301 VGND.n924 VGND.n836 2306.06
R302 VGND.n924 VGND.n840 2306.06
R303 VGND.n930 VGND.n825 2306.06
R304 VGND.n825 VGND.n780 2306.06
R305 VGND.n896 VGND.n892 2306.06
R306 VGND.n896 VGND.n893 2306.06
R307 VGND.n915 VGND.n842 2306.06
R308 VGND.n915 VGND.n843 2306.06
R309 VGND.n886 VGND.n861 2306.06
R310 VGND.n890 VGND.n861 2306.06
R311 VGND.n886 VGND.n862 2306.06
R312 VGND.n890 VGND.n862 2306.06
R313 VGND.n873 VGND.n872 2306.06
R314 VGND.n872 VGND.n864 2306.06
R315 VGND.n874 VGND.n873 2306.06
R316 VGND.n874 VGND.n864 2306.06
R317 VGND.n969 VGND.n261 2306.06
R318 VGND.n973 VGND.n261 2306.06
R319 VGND.n969 VGND.n262 2306.06
R320 VGND.n973 VGND.n262 2306.06
R321 VGND.n803 VGND.n265 2168.06
R322 VGND.n1025 VGND.n1024 2024.56
R323 VGND.n672 VGND.n450 1455.1
R324 VGND.n689 VGND.n454 1455.1
R325 VGND.n731 VGND.n281 1455.1
R326 VGND.n749 VGND.n284 1455.1
R327 VGND.n124 VGND.n34 1455.1
R328 VGND.n1003 VGND.n37 1455.1
R329 VGND.n1022 VGND.n15 1401.31
R330 VGND.n510 VGND.n509 1390.59
R331 VGND.n509 VGND.n505 1390.59
R332 VGND.n511 VGND.n508 1390.59
R333 VGND.n511 VGND.n504 1390.59
R334 VGND.n775 VGND.n771 1390.59
R335 VGND.n775 VGND.n765 1390.59
R336 VGND.n772 VGND.n770 1390.59
R337 VGND.n772 VGND.n764 1390.59
R338 VGND.n828 VGND.n824 1390.59
R339 VGND.n828 VGND.n827 1390.59
R340 VGND.n838 VGND.n837 1390.59
R341 VGND.n839 VGND.n838 1390.59
R342 VGND.n852 VGND.n851 1390.59
R343 VGND.n851 VGND.n847 1390.59
R344 VGND.n853 VGND.n850 1390.59
R345 VGND.n853 VGND.n846 1390.59
R346 VGND.n672 VGND.n473 1389.8
R347 VGND.n689 VGND.n450 1389.8
R348 VGND.n731 VGND.n407 1389.8
R349 VGND.n749 VGND.n281 1389.8
R350 VGND.n124 VGND.n66 1389.8
R351 VGND.n1003 VGND.n34 1389.8
R352 VGND.n161 VGND.n150 1373.21
R353 VGND.n165 VGND.n164 1373.21
R354 VGND.n164 VGND.n148 1373.21
R355 VGND.n156 VGND.n148 1373.21
R356 VGND.n169 VGND.n139 1373.21
R357 VGND.n169 VGND.n142 1373.21
R358 VGND.n162 VGND.n142 1373.21
R359 VGND.n162 VGND.n161 1373.21
R360 VGND.n139 VGND.n137 1373.21
R361 VGND.n174 VGND.n173 1373.21
R362 VGND.n173 VGND.n138 1373.21
R363 VGND.n165 VGND.n138 1373.21
R364 VGND.n954 VGND.n953 1320.82
R365 VGND.n965 VGND.n954 1320.82
R366 VGND.n186 VGND.n182 1309.47
R367 VGND.n191 VGND.n188 1309.47
R368 VGND.n191 VGND.n7 1309.47
R369 VGND.n195 VGND.n8 1309.47
R370 VGND.n214 VGND.n213 1309.47
R371 VGND.n214 VGND.n195 1309.47
R372 VGND.n210 VGND.n199 1309.47
R373 VGND.n199 VGND.n188 1309.47
R374 VGND.n203 VGND.n200 1309.47
R375 VGND.n203 VGND.n186 1309.47
R376 VGND.n81 VGND.n63 1309.47
R377 VGND.n67 VGND.n65 1309.47
R378 VGND.n68 VGND.n67 1309.47
R379 VGND.n997 VGND.n45 1309.47
R380 VGND.n998 VGND.n41 1309.47
R381 VGND.n998 VGND.n997 1309.47
R382 VGND.n64 VGND.n40 1309.47
R383 VGND.n65 VGND.n64 1309.47
R384 VGND.n74 VGND.n73 1309.47
R385 VGND.n74 VGND.n63 1309.47
R386 VGND.n102 VGND.n32 1309.47
R387 VGND.n103 VGND.n102 1309.47
R388 VGND.n91 VGND.n88 1309.47
R389 VGND.n107 VGND.n33 1309.47
R390 VGND.n94 VGND.n88 1309.47
R391 VGND.n94 VGND.n93 1309.47
R392 VGND.n105 VGND.n103 1309.47
R393 VGND.n105 VGND.n104 1309.47
R394 VGND.n108 VGND.n107 1309.47
R395 VGND.n108 VGND.n54 1309.47
R396 VGND.n435 VGND.n434 1309.47
R397 VGND.n705 VGND.n703 1309.47
R398 VGND.n705 VGND.n704 1309.47
R399 VGND.n743 VGND.n292 1309.47
R400 VGND.n744 VGND.n288 1309.47
R401 VGND.n744 VGND.n743 1309.47
R402 VGND.n702 VGND.n287 1309.47
R403 VGND.n703 VGND.n702 1309.47
R404 VGND.n433 VGND.n412 1309.47
R405 VGND.n434 VGND.n433 1309.47
R406 VGND.n637 VGND.n636 1309.47
R407 VGND.n641 VGND.n448 1309.47
R408 VGND.n641 VGND.n640 1309.47
R409 VGND.n645 VGND.n449 1309.47
R410 VGND.n684 VGND.n457 1309.47
R411 VGND.n684 VGND.n449 1309.47
R412 VGND.n458 VGND.n456 1309.47
R413 VGND.n458 VGND.n448 1309.47
R414 VGND.n635 VGND.n478 1309.47
R415 VGND.n636 VGND.n635 1309.47
R416 VGND.n424 VGND.n423 1309.47
R417 VGND.n424 VGND.n279 1309.47
R418 VGND.n716 VGND.n420 1309.47
R419 VGND.n427 VGND.n280 1309.47
R420 VGND.n718 VGND.n420 1309.47
R421 VGND.n718 VGND.n404 1309.47
R422 VGND.n405 VGND.n279 1309.47
R423 VGND.n406 VGND.n405 1309.47
R424 VGND.n400 VGND.n280 1309.47
R425 VGND.n400 VGND.n398 1309.47
R426 VGND.n624 VGND.n621 1309.47
R427 VGND.n624 VGND.n623 1309.47
R428 VGND.n616 VGND.n613 1309.47
R429 VGND.n655 VGND.n654 1309.47
R430 VGND.n618 VGND.n613 1309.47
R431 VGND.n618 VGND.n471 1309.47
R432 VGND.n623 VGND.n622 1309.47
R433 VGND.n622 VGND.n472 1309.47
R434 VGND.n654 VGND.n653 1309.47
R435 VGND.n653 VGND.n466 1309.47
R436 VGND.n666 VGND.n609 1136.73
R437 VGND.n666 VGND.n473 1136.73
R438 VGND.n681 VGND.n454 1136.73
R439 VGND.n681 VGND.n465 1136.73
R440 VGND.n725 VGND.n416 1136.73
R441 VGND.n725 VGND.n407 1136.73
R442 VGND.n741 VGND.n284 1136.73
R443 VGND.n741 VGND.n397 1136.73
R444 VGND.n118 VGND.n78 1136.73
R445 VGND.n118 VGND.n66 1136.73
R446 VGND.n995 VGND.n37 1136.73
R447 VGND.n995 VGND.n53 1136.73
R448 VGND.n965 VGND.n964 1057.25
R449 VGND.n547 VGND.n508 915.471
R450 VGND.n552 VGND.n508 915.471
R451 VGND.n552 VGND.n510 915.471
R452 VGND.n510 VGND.n499 915.471
R453 VGND.n545 VGND.n504 915.471
R454 VGND.n554 VGND.n504 915.471
R455 VGND.n554 VGND.n505 915.471
R456 VGND.n505 VGND.n500 915.471
R457 VGND.n918 VGND.n770 915.471
R458 VGND.n936 VGND.n770 915.471
R459 VGND.n936 VGND.n771 915.471
R460 VGND.n932 VGND.n771 915.471
R461 VGND.n919 VGND.n764 915.471
R462 VGND.n938 VGND.n764 915.471
R463 VGND.n938 VGND.n765 915.471
R464 VGND.n779 VGND.n765 915.471
R465 VGND.n837 VGND.n836 915.471
R466 VGND.n837 VGND.n769 915.471
R467 VGND.n824 VGND.n769 915.471
R468 VGND.n930 VGND.n824 915.471
R469 VGND.n840 VGND.n839 915.471
R470 VGND.n839 VGND.n767 915.471
R471 VGND.n827 VGND.n767 915.471
R472 VGND.n827 VGND.n780 915.471
R473 VGND.n892 VGND.n850 915.471
R474 VGND.n908 VGND.n850 915.471
R475 VGND.n908 VGND.n852 915.471
R476 VGND.n852 VGND.n842 915.471
R477 VGND.n893 VGND.n846 915.471
R478 VGND.n910 VGND.n846 915.471
R479 VGND.n910 VGND.n847 915.471
R480 VGND.n847 VGND.n843 915.471
R481 VGND.n465 VGND.n416 751.02
R482 VGND.n180 VGND.n53 751.02
R483 VGND.n1024 VGND.n1023 727.957
R484 VGND.n243 VGND.n242 705.365
R485 VGND.n350 VGND.n347 666.73
R486 VGND VGND.n350 666.73
R487 VGND.n1021 VGND.n1020 665.898
R488 VGND.n235 VGND.n180 659.184
R489 VGND.n949 VGND.n269 621.553
R490 VGND.n948 VGND 619.196
R491 VGND.n242 VGND.n241 599.019
R492 VGND.n951 VGND.n266 578.904
R493 VGND.n308 VGND.n266 578.904
R494 VGND.n315 VGND.n308 578.904
R495 VGND.n315 VGND.n296 578.904
R496 VGND.n395 VGND.n298 578.904
R497 VGND.n387 VGND.n298 578.904
R498 VGND.n387 VGND.n320 578.904
R499 VGND.n383 VGND.n320 578.904
R500 VGND.n383 VGND.n382 578.904
R501 VGND.n382 VGND.n325 578.904
R502 VGND.n375 VGND.n325 578.904
R503 VGND.n375 VGND.n374 578.904
R504 VGND.n374 VGND.n335 578.904
R505 VGND.n366 VGND.n335 578.904
R506 VGND.n366 VGND.n343 578.904
R507 VGND.n343 VGND.n12 578.904
R508 VGND.n353 VGND.n13 578.904
R509 VGND.n353 VGND.n351 578.904
R510 VGND.n524 VGND.n263 560.645
R511 VGND.n528 VGND.n524 560.645
R512 VGND.n527 VGND.n515 560.645
R513 VGND.n542 VGND.n515 560.645
R514 VGND.n546 VGND.n543 560.645
R515 VGND.n546 VGND.n506 560.645
R516 VGND.n553 VGND.n506 560.645
R517 VGND.n553 VGND.n507 560.645
R518 VGND.n507 VGND.n498 560.645
R519 VGND.n558 VGND.n498 560.645
R520 VGND.n561 VGND.n489 560.645
R521 VGND.n571 VGND.n489 560.645
R522 VGND.n574 VGND.n482 560.645
R523 VGND.n585 VGND.n482 560.645
R524 VGND.n863 VGND.n264 560.645
R525 VGND.n882 VGND.n863 560.645
R526 VGND.n885 VGND.n860 560.645
R527 VGND.n898 VGND.n860 560.645
R528 VGND.n897 VGND.n891 560.645
R529 VGND.n891 VGND.n848 560.645
R530 VGND.n909 VGND.n848 560.645
R531 VGND.n909 VGND.n849 560.645
R532 VGND.n849 VGND.n841 560.645
R533 VGND.n916 VGND.n841 560.645
R534 VGND.n923 VGND.n917 560.645
R535 VGND.n917 VGND.n766 560.645
R536 VGND.n937 VGND.n766 560.645
R537 VGND.n937 VGND.n768 560.645
R538 VGND.n931 VGND.n768 560.645
R539 VGND.n931 VGND.n823 560.645
R540 VGND.n822 VGND.n782 560.645
R541 VGND.n814 VGND.n782 560.645
R542 VGND.n812 VGND.n792 560.645
R543 VGND.n803 VGND.n792 560.645
R544 VGND.n968 VGND.n259 560.645
R545 VGND.n974 VGND.n259 560.645
R546 VGND.n586 VGND.n260 560.645
R547 VGND.n605 VGND.n586 560.645
R548 VGND.n152 VGND 551.907
R549 VGND.n157 VGND.n152 551.907
R550 VGND.n176 VGND.n136 551.907
R551 VGND.n237 VGND.n235 550.859
R552 VGND.n1023 VGND.n13 530.803
R553 VGND.n211 VGND.n196 490.01
R554 VGND.n221 VGND.n196 490.01
R555 VGND.n221 VGND.n9 490.01
R556 VGND.n1025 VGND.n9 490.01
R557 VGND.n159 VGND.n151 462.683
R558 VGND.n159 VGND.n158 462.683
R559 VGND.n168 VGND.n167 462.683
R560 VGND.n167 VGND.n147 462.683
R561 VGND.n143 VGND.n140 462.683
R562 VGND.n145 VGND.n140 462.683
R563 VGND.n171 VGND.n11 435.882
R564 VGND.n171 VGND.n170 435.882
R565 VGND.n170 VGND.n141 435.882
R566 VGND.n163 VGND.n141 435.882
R567 VGND.n163 VGND.n149 435.882
R568 VGND.n155 VGND.n149 435.882
R569 VGND.n154 VGND.n153 424.591
R570 VGND.n208 VGND.n187 417.005
R571 VGND.n227 VGND.n187 417.005
R572 VGND.n227 VGND.n181 417.005
R573 VGND.n234 VGND.n181 417.005
R574 VGND.n238 VGND.n237 417.005
R575 VGND.n239 VGND.n238 417.005
R576 VGND.n361 VGND.n360 414.872
R577 VGND.n360 VGND.n348 414.872
R578 VGND.n355 VGND.n346 414.872
R579 VGND.n356 VGND.n355 414.872
R580 VGND.n339 VGND.n334 414.872
R581 VGND.n334 VGND.n331 414.872
R582 VGND.n371 VGND.n370 414.872
R583 VGND.n370 VGND.n341 414.872
R584 VGND.n380 VGND.n327 414.872
R585 VGND.n380 VGND.n379 414.872
R586 VGND.n329 VGND.n328 414.872
R587 VGND.n330 VGND.n329 414.872
R588 VGND.n303 VGND.n301 414.872
R589 VGND.n317 VGND.n303 414.872
R590 VGND.n392 VGND.n391 414.872
R591 VGND.n391 VGND.n318 414.872
R592 VGND.n312 VGND.n311 414.872
R593 VGND.n311 VGND.n304 414.872
R594 VGND.n561 VGND.n558 376.13
R595 VGND.n898 VGND.n897 376.13
R596 VGND.n923 VGND.n916 376.13
R597 VGND.n823 VGND.n822 376.13
R598 VGND.n528 VGND.n527 369.033
R599 VGND.n574 VGND.n571 369.033
R600 VGND.n885 VGND.n882 369.033
R601 VGND.n814 VGND.n812 369.033
R602 VGND.n974 VGND.n260 369.033
R603 VGND.n396 VGND.n395 360.339
R604 VGND.n926 VGND.n925 343.154
R605 VGND.n1024 VGND.n11 339.783
R606 VGND.n177 VGND 335.06
R607 VGND.n97 VGND.n89 294.776
R608 VGND.n615 VGND.n614 294.776
R609 VGND.n293 VGND.n290 294.776
R610 VGND.n422 VGND.n421 294.776
R611 VGND.n738 VGND.n737 294.776
R612 VGND.n727 VGND.n414 294.776
R613 VGND.n683 VGND.n461 294.776
R614 VGND.n668 VGND.n480 294.776
R615 VGND.n679 VGND.n678 294.776
R616 VGND.n218 VGND.n217 294.776
R617 VGND.n206 VGND.n184 294.776
R618 VGND.n50 VGND.n43 294.776
R619 VGND.n120 VGND.n76 294.776
R620 VGND.n992 VGND.n991 294.776
R621 VGND.n564 VGND.n563 292.5
R622 VGND.n563 VGND.n489 292.5
R623 VGND.n497 VGND 292.5
R624 VGND.n497 VGND.n489 292.5
R625 VGND.n577 VGND.n576 292.5
R626 VGND.n576 VGND.n482 292.5
R627 VGND.n488 VGND 292.5
R628 VGND.n488 VGND.n482 292.5
R629 VGND.n523 VGND 292.5
R630 VGND.n524 VGND.n523 292.5
R631 VGND.n520 VGND.n519 292.5
R632 VGND.n524 VGND.n520 292.5
R633 VGND VGND.n517 292.5
R634 VGND.n517 VGND.n515 292.5
R635 VGND.n518 VGND.n516 292.5
R636 VGND.n516 VGND.n515 292.5
R637 VGND VGND.n500 292.5
R638 VGND.n500 VGND.n498 292.5
R639 VGND VGND.n554 292.5
R640 VGND.n554 VGND.n553 292.5
R641 VGND.n545 VGND 292.5
R642 VGND.n546 VGND.n545 292.5
R643 VGND.n548 VGND.n547 292.5
R644 VGND.n547 VGND.n546 292.5
R645 VGND.n552 VGND.n551 292.5
R646 VGND.n553 VGND.n552 292.5
R647 VGND.n501 VGND.n499 292.5
R648 VGND.n499 VGND.n498 292.5
R649 VGND VGND.n492 292.5
R650 VGND.n492 VGND.n489 292.5
R651 VGND.n493 VGND.n491 292.5
R652 VGND.n491 VGND.n489 292.5
R653 VGND VGND.n485 292.5
R654 VGND.n485 VGND.n482 292.5
R655 VGND.n486 VGND.n484 292.5
R656 VGND.n484 VGND.n482 292.5
R657 VGND.n875 VGND.n874 292.5
R658 VGND.n874 VGND.n863 292.5
R659 VGND.n872 VGND 292.5
R660 VGND.n872 VGND.n863 292.5
R661 VGND.n888 VGND.n862 292.5
R662 VGND.n862 VGND.n860 292.5
R663 VGND VGND.n861 292.5
R664 VGND.n861 VGND.n860 292.5
R665 VGND.n913 VGND.n843 292.5
R666 VGND.n843 VGND.n841 292.5
R667 VGND.n911 VGND.n910 292.5
R668 VGND.n910 VGND.n909 292.5
R669 VGND.n894 VGND.n893 292.5
R670 VGND.n893 VGND.n891 292.5
R671 VGND VGND.n892 292.5
R672 VGND.n892 VGND.n891 292.5
R673 VGND.n908 VGND 292.5
R674 VGND.n909 VGND.n908 292.5
R675 VGND VGND.n842 292.5
R676 VGND.n842 VGND.n841 292.5
R677 VGND.n831 VGND.n780 292.5
R678 VGND.n931 VGND.n780 292.5
R679 VGND.n833 VGND.n767 292.5
R680 VGND.n937 VGND.n767 292.5
R681 VGND.n840 VGND.n835 292.5
R682 VGND.n917 VGND.n840 292.5
R683 VGND.n836 VGND 292.5
R684 VGND.n917 VGND.n836 292.5
R685 VGND VGND.n769 292.5
R686 VGND.n937 VGND.n769 292.5
R687 VGND.n930 VGND 292.5
R688 VGND.n931 VGND.n930 292.5
R689 VGND.n790 VGND.n788 292.5
R690 VGND.n790 VGND.n782 292.5
R691 VGND.n789 VGND 292.5
R692 VGND.n789 VGND.n782 292.5
R693 VGND.n801 VGND.n799 292.5
R694 VGND.n801 VGND.n792 292.5
R695 VGND.n800 VGND 292.5
R696 VGND.n800 VGND.n792 292.5
R697 VGND VGND.n866 292.5
R698 VGND.n866 VGND.n863 292.5
R699 VGND.n867 VGND.n865 292.5
R700 VGND.n865 VGND.n863 292.5
R701 VGND.n859 VGND 292.5
R702 VGND.n860 VGND.n859 292.5
R703 VGND.n858 VGND.n857 292.5
R704 VGND.n860 VGND.n858 292.5
R705 VGND.n779 VGND 292.5
R706 VGND.n931 VGND.n779 292.5
R707 VGND VGND.n938 292.5
R708 VGND.n938 VGND.n937 292.5
R709 VGND VGND.n919 292.5
R710 VGND.n919 VGND.n917 292.5
R711 VGND.n920 VGND.n918 292.5
R712 VGND.n918 VGND.n917 292.5
R713 VGND.n936 VGND.n935 292.5
R714 VGND.n937 VGND.n936 292.5
R715 VGND.n933 VGND.n932 292.5
R716 VGND.n932 VGND.n931 292.5
R717 VGND VGND.n784 292.5
R718 VGND.n784 VGND.n782 292.5
R719 VGND.n785 VGND.n783 292.5
R720 VGND.n783 VGND.n782 292.5
R721 VGND VGND.n794 292.5
R722 VGND.n794 VGND.n792 292.5
R723 VGND.n795 VGND.n793 292.5
R724 VGND.n793 VGND.n792 292.5
R725 VGND VGND.n18 292.5
R726 VGND.n1020 VGND.n18 292.5
R727 VGND.n961 VGND.n960 292.5
R728 VGND.n964 VGND.n961 292.5
R729 VGND.n1019 VGND 292.5
R730 VGND.n1020 VGND.n1019 292.5
R731 VGND.n963 VGND.n962 292.5
R732 VGND.n964 VGND.n963 292.5
R733 VGND.n597 VGND.n596 292.5
R734 VGND.n596 VGND.n586 292.5
R735 VGND.n594 VGND 292.5
R736 VGND.n594 VGND.n586 292.5
R737 VGND.n258 VGND 292.5
R738 VGND.n259 VGND.n258 292.5
R739 VGND.n257 VGND.n256 292.5
R740 VGND.n259 VGND.n257 292.5
R741 VGND VGND.n589 292.5
R742 VGND.n589 VGND.n586 292.5
R743 VGND.n590 VGND.n588 292.5
R744 VGND.n588 VGND.n586 292.5
R745 VGND.n971 VGND.n262 292.5
R746 VGND.n262 VGND.n259 292.5
R747 VGND VGND.n261 292.5
R748 VGND.n261 VGND.n259 292.5
R749 VGND VGND.n178 289.281
R750 VGND VGND.n134 285.604
R751 VGND.n429 VGND.n428 280.32
R752 VGND.n710 VGND.n709 280.32
R753 VGND.n647 VGND.n646 280.32
R754 VGND.n656 VGND.n652 280.32
R755 VGND.n1027 VGND.n6 280.32
R756 VGND.n48 VGND.n47 280.32
R757 VGND.n1005 VGND.n31 280.32
R758 VGND.n734 VGND.n733 268.425
R759 VGND.n736 VGND.n735 268.425
R760 VGND.n715 VGND.n714 268.425
R761 VGND.n707 VGND.n432 268.425
R762 VGND.n729 VGND.n289 268.425
R763 VGND.n747 VGND.n746 268.425
R764 VGND.n643 VGND.n639 268.425
R765 VGND.n670 VGND.n460 268.425
R766 VGND.n687 VGND.n686 268.425
R767 VGND.n627 VGND.n626 268.425
R768 VGND.n675 VGND.n674 268.425
R769 VGND.n677 VGND.n676 268.425
R770 VGND.n232 VGND.n5 268.425
R771 VGND.n202 VGND.n201 268.425
R772 VGND.n216 VGND.n198 268.425
R773 VGND.n80 VGND.n79 268.425
R774 VGND.n122 VGND.n42 268.425
R775 VGND.n1001 VGND.n1000 268.425
R776 VGND.n90 VGND.n30 268.425
R777 VGND.n101 VGND.n99 268.425
R778 VGND.n100 VGND.n56 268.425
R779 VGND.n717 VGND.n715 268.274
R780 VGND.n436 VGND.n432 268.274
R781 VGND.n639 VGND.n638 268.274
R782 VGND.n626 VGND.n617 268.274
R783 VGND.n232 VGND.n231 268.274
R784 VGND.n82 VGND.n80 268.274
R785 VGND.n92 VGND.n90 268.274
R786 VGND.n733 VGND.n403 256.377
R787 VGND.n735 VGND.n734 256.377
R788 VGND.n729 VGND.n728 256.377
R789 VGND.n747 VGND.n289 256.377
R790 VGND.n670 VGND.n669 256.377
R791 VGND.n687 VGND.n460 256.377
R792 VGND.n674 VGND.n470 256.377
R793 VGND.n676 VGND.n675 256.377
R794 VGND.n205 VGND.n202 256.377
R795 VGND.n201 VGND.n198 256.377
R796 VGND.n122 VGND.n121 256.377
R797 VGND.n1001 VGND.n42 256.377
R798 VGND.n99 VGND.n98 256.377
R799 VGND.n101 VGND.n100 256.377
R800 VGND.n713 VGND.n429 256
R801 VGND.n711 VGND.n710 256
R802 VGND.n648 VGND.n647 256
R803 VGND.n652 VGND.n651 256
R804 VGND.n1028 VGND.n1027 256
R805 VGND.n47 VGND.n28 256
R806 VGND.n1006 VGND.n1005 256
R807 VGND.n313 VGND.n312 251.859
R808 VGND.n313 VGND.n301 251.859
R809 VGND.n338 VGND.n327 251.859
R810 VGND.n339 VGND.n338 251.859
R811 VGND.n361 VGND.n347 251.859
R812 VGND VGND.n356 251.859
R813 VGND VGND.n348 251.859
R814 VGND VGND.n348 251.859
R815 VGND.n371 VGND.n340 251.859
R816 VGND.n346 VGND.n340 251.859
R817 VGND.n362 VGND.n346 251.859
R818 VGND.n362 VGND.n361 251.859
R819 VGND VGND.n331 251.859
R820 VGND.n341 VGND 251.859
R821 VGND VGND.n341 251.859
R822 VGND.n356 VGND 251.859
R823 VGND.n372 VGND.n339 251.859
R824 VGND.n372 VGND.n371 251.859
R825 VGND VGND.n330 251.859
R826 VGND.n379 VGND 251.859
R827 VGND.n379 VGND 251.859
R828 VGND VGND.n331 251.859
R829 VGND.n392 VGND.n302 251.859
R830 VGND.n328 VGND.n302 251.859
R831 VGND.n328 VGND.n323 251.859
R832 VGND.n327 VGND.n323 251.859
R833 VGND VGND.n317 251.859
R834 VGND.n318 VGND 251.859
R835 VGND VGND.n318 251.859
R836 VGND.n330 VGND 251.859
R837 VGND.n393 VGND.n301 251.859
R838 VGND.n393 VGND.n392 251.859
R839 VGND.n304 VGND 251.859
R840 VGND VGND.n304 251.859
R841 VGND.n317 VGND 251.859
R842 VGND.n312 VGND.n269 251.859
R843 VGND.n929 VGND.n928 249.667
R844 VGND.n396 VGND.n296 218.565
R845 VGND.n177 VGND.n176 216.847
R846 VGND.n421 VGND.n403 209.695
R847 VGND.n738 VGND.n736 209.695
R848 VGND.n728 VGND.n727 209.695
R849 VGND.n746 VGND.n290 209.695
R850 VGND.n669 VGND.n668 209.695
R851 VGND.n686 VGND.n683 209.695
R852 VGND.n614 VGND.n470 209.695
R853 VGND.n679 VGND.n677 209.695
R854 VGND.n206 VGND.n205 209.695
R855 VGND.n217 VGND.n216 209.695
R856 VGND.n121 VGND.n120 209.695
R857 VGND.n1000 VGND.n43 209.695
R858 VGND.n98 VGND.n97 209.695
R859 VGND.n992 VGND.n56 209.695
R860 VGND.n954 VGND.n263 188.065
R861 VGND.n607 VGND.n585 188.065
R862 VGND.n953 VGND.n264 188.065
R863 VGND.n606 VGND.n605 188.065
R864 VGND.n239 VGND.n10 151.014
R865 VGND.n556 VGND.n501 150.417
R866 VGND.n933 VGND.n777 150.417
R867 VGND.n831 VGND.n826 150.417
R868 VGND.n914 VGND.n913 150.417
R869 VGND.n592 VGND.n590 149.835
R870 VGND.n603 VGND.n590 149.835
R871 VGND VGND.n592 149.835
R872 VGND.n966 VGND.n256 149.835
R873 VGND.n976 VGND.n256 149.835
R874 VGND.n966 VGND 149.835
R875 VGND.n593 VGND 149.835
R876 VGND.n597 VGND.n593 149.835
R877 VGND.n598 VGND.n597 149.835
R878 VGND.n572 VGND.n486 149.835
R879 VGND.n572 VGND 149.835
R880 VGND.n583 VGND.n486 149.835
R881 VGND.n559 VGND.n493 149.835
R882 VGND.n559 VGND 149.835
R883 VGND.n569 VGND.n493 149.835
R884 VGND.n548 VGND.n513 149.835
R885 VGND.n525 VGND.n518 149.835
R886 VGND.n525 VGND 149.835
R887 VGND.n540 VGND.n518 149.835
R888 VGND.n521 VGND.n519 149.835
R889 VGND.n521 VGND 149.835
R890 VGND.n530 VGND.n519 149.835
R891 VGND.n578 VGND.n577 149.835
R892 VGND.n577 VGND.n487 149.835
R893 VGND.n487 VGND 149.835
R894 VGND.n496 VGND 149.835
R895 VGND.n564 VGND.n496 149.835
R896 VGND.n565 VGND.n564 149.835
R897 VGND.n810 VGND.n795 149.835
R898 VGND.n810 VGND 149.835
R899 VGND.n796 VGND.n795 149.835
R900 VGND.n820 VGND.n785 149.835
R901 VGND.n820 VGND 149.835
R902 VGND.n786 VGND.n785 149.835
R903 VGND.n921 VGND.n920 149.835
R904 VGND.n883 VGND.n857 149.835
R905 VGND.n883 VGND 149.835
R906 VGND.n900 VGND.n857 149.835
R907 VGND.n869 VGND.n867 149.835
R908 VGND VGND.n869 149.835
R909 VGND.n880 VGND.n867 149.835
R910 VGND.n805 VGND.n799 149.835
R911 VGND.n799 VGND.n798 149.835
R912 VGND.n798 VGND 149.835
R913 VGND.n816 VGND.n788 149.835
R914 VGND.n788 VGND.n787 149.835
R915 VGND.n787 VGND 149.835
R916 VGND.n889 VGND.n888 149.835
R917 VGND.n888 VGND.n887 149.835
R918 VGND.n887 VGND 149.835
R919 VGND.n925 VGND.n835 149.835
R920 VGND.n895 VGND.n894 149.835
R921 VGND.n871 VGND 149.835
R922 VGND.n875 VGND.n871 149.835
R923 VGND.n876 VGND.n875 149.835
R924 VGND.n962 VGND.n21 149.835
R925 VGND VGND.n21 149.835
R926 VGND.n962 VGND.n22 149.835
R927 VGND.n960 VGND.n957 149.835
R928 VGND VGND.n957 149.835
R929 VGND.n960 VGND.n959 149.835
R930 VGND.n972 VGND.n971 149.835
R931 VGND.n971 VGND.n970 149.835
R932 VGND.n970 VGND 149.835
R933 VGND.n603 VGND.n602 149.459
R934 VGND.n977 VGND.n976 149.459
R935 VGND.n599 VGND.n598 149.459
R936 VGND.n583 VGND.n582 149.459
R937 VGND.n569 VGND.n568 149.459
R938 VGND.n540 VGND.n539 149.459
R939 VGND.n531 VGND.n530 149.459
R940 VGND.n579 VGND.n578 149.459
R941 VGND.n566 VGND.n565 149.459
R942 VGND.n809 VGND.n796 149.459
R943 VGND.n819 VGND.n786 149.459
R944 VGND.n901 VGND.n900 149.459
R945 VGND.n880 VGND.n879 149.459
R946 VGND.n806 VGND.n805 149.459
R947 VGND.n817 VGND.n816 149.459
R948 VGND.n889 VGND.n856 149.459
R949 VGND.n877 VGND.n876 149.459
R950 VGND.n1018 VGND.n22 149.459
R951 VGND.n959 VGND.n958 149.459
R952 VGND.n972 VGND.n255 149.459
R953 VGND.n928 VGND.n927 132.8
R954 VGND.n914 VGND 132.129
R955 VGND.n556 VGND 132.127
R956 VGND VGND.n777 132.127
R957 VGND VGND.n513 130.802
R958 VGND.n921 VGND 130.802
R959 VGND.n895 VGND 130.802
R960 VGND VGND.n178 130.327
R961 VGND.n927 VGND.n926 120.001
R962 VGND VGND 118.966
R963 VGND.n242 VGND.n135 117.272
R964 VGND.n565 VGND.n490 117.001
R965 VGND.n571 VGND.n490 117.001
R966 VGND.n562 VGND.n496 117.001
R967 VGND.n562 VGND.n561 117.001
R968 VGND.n578 VGND.n483 117.001
R969 VGND.n585 VGND.n483 117.001
R970 VGND.n575 VGND.n487 117.001
R971 VGND.n575 VGND.n574 117.001
R972 VGND.n530 VGND.n529 117.001
R973 VGND.n529 VGND.n528 117.001
R974 VGND.n522 VGND.n521 117.001
R975 VGND.n522 VGND.n263 117.001
R976 VGND.n541 VGND.n540 117.001
R977 VGND.n542 VGND.n541 117.001
R978 VGND.n526 VGND.n525 117.001
R979 VGND.n527 VGND.n526 117.001
R980 VGND.n512 VGND.n511 117.001
R981 VGND.n511 VGND.n506 117.001
R982 VGND.n509 VGND.n502 117.001
R983 VGND.n509 VGND.n507 117.001
R984 VGND.n557 VGND.n556 117.001
R985 VGND.n558 VGND.n557 117.001
R986 VGND.n514 VGND.n513 117.001
R987 VGND.n543 VGND.n514 117.001
R988 VGND.n570 VGND.n569 117.001
R989 VGND.n571 VGND.n570 117.001
R990 VGND.n560 VGND.n559 117.001
R991 VGND.n561 VGND.n560 117.001
R992 VGND.n584 VGND.n583 117.001
R993 VGND.n585 VGND.n584 117.001
R994 VGND.n573 VGND.n572 117.001
R995 VGND.n574 VGND.n573 117.001
R996 VGND.n876 VGND.n864 117.001
R997 VGND.n882 VGND.n864 117.001
R998 VGND.n873 VGND.n871 117.001
R999 VGND.n873 VGND.n264 117.001
R1000 VGND.n890 VGND.n889 117.001
R1001 VGND.n898 VGND.n890 117.001
R1002 VGND.n887 VGND.n886 117.001
R1003 VGND.n886 VGND.n885 117.001
R1004 VGND.n854 VGND.n853 117.001
R1005 VGND.n853 VGND.n848 117.001
R1006 VGND.n851 VGND.n844 117.001
R1007 VGND.n851 VGND.n849 117.001
R1008 VGND.n915 VGND.n914 117.001
R1009 VGND.n916 VGND.n915 117.001
R1010 VGND.n896 VGND.n895 117.001
R1011 VGND.n897 VGND.n896 117.001
R1012 VGND.n838 VGND.n830 117.001
R1013 VGND.n838 VGND.n766 117.001
R1014 VGND.n829 VGND.n828 117.001
R1015 VGND.n828 VGND.n768 117.001
R1016 VGND.n826 VGND.n825 117.001
R1017 VGND.n825 VGND.n823 117.001
R1018 VGND.n925 VGND.n924 117.001
R1019 VGND.n924 VGND.n923 117.001
R1020 VGND.n816 VGND.n815 117.001
R1021 VGND.n815 VGND.n814 117.001
R1022 VGND.n787 VGND.n781 117.001
R1023 VGND.n822 VGND.n781 117.001
R1024 VGND.n805 VGND.n804 117.001
R1025 VGND.n804 VGND.n803 117.001
R1026 VGND.n798 VGND.n791 117.001
R1027 VGND.n812 VGND.n791 117.001
R1028 VGND.n881 VGND.n880 117.001
R1029 VGND.n882 VGND.n881 117.001
R1030 VGND.n869 VGND.n868 117.001
R1031 VGND.n868 VGND.n264 117.001
R1032 VGND.n900 VGND.n899 117.001
R1033 VGND.n899 VGND.n898 117.001
R1034 VGND.n884 VGND.n883 117.001
R1035 VGND.n885 VGND.n884 117.001
R1036 VGND.n773 VGND.n772 117.001
R1037 VGND.n772 VGND.n766 117.001
R1038 VGND.n776 VGND.n775 117.001
R1039 VGND.n775 VGND.n768 117.001
R1040 VGND.n778 VGND.n777 117.001
R1041 VGND.n823 VGND.n778 117.001
R1042 VGND.n922 VGND.n921 117.001
R1043 VGND.n923 VGND.n922 117.001
R1044 VGND.n813 VGND.n786 117.001
R1045 VGND.n814 VGND.n813 117.001
R1046 VGND.n821 VGND.n820 117.001
R1047 VGND.n822 VGND.n821 117.001
R1048 VGND.n802 VGND.n796 117.001
R1049 VGND.n803 VGND.n802 117.001
R1050 VGND.n811 VGND.n810 117.001
R1051 VGND.n812 VGND.n811 117.001
R1052 VGND.n619 VGND.n618 117.001
R1053 VGND.n618 VGND.n473 117.001
R1054 VGND.n656 VGND.n655 117.001
R1055 VGND.n655 VGND.n454 117.001
R1056 VGND.n653 VGND.n468 117.001
R1057 VGND.n653 VGND.n454 117.001
R1058 VGND.n625 VGND.n624 117.001
R1059 VGND.n624 VGND.n450 117.001
R1060 VGND.n622 VGND.n469 117.001
R1061 VGND.n622 VGND.n450 117.001
R1062 VGND.n678 VGND.n467 117.001
R1063 VGND.n467 VGND.n465 117.001
R1064 VGND.n615 VGND.n612 117.001
R1065 VGND.n612 VGND.n609 117.001
R1066 VGND.n617 VGND.n616 117.001
R1067 VGND.n616 VGND.n473 117.001
R1068 VGND.n719 VGND.n718 117.001
R1069 VGND.n718 VGND.n407 117.001
R1070 VGND.n428 VGND.n427 117.001
R1071 VGND.n427 VGND.n284 117.001
R1072 VGND.n401 VGND.n400 117.001
R1073 VGND.n400 VGND.n284 117.001
R1074 VGND.n425 VGND.n424 117.001
R1075 VGND.n424 VGND.n281 117.001
R1076 VGND.n405 VGND.n402 117.001
R1077 VGND.n405 VGND.n281 117.001
R1078 VGND.n737 VGND.n399 117.001
R1079 VGND.n399 VGND.n397 117.001
R1080 VGND.n422 VGND.n419 117.001
R1081 VGND.n419 VGND.n416 117.001
R1082 VGND.n717 VGND.n716 117.001
R1083 VGND.n716 VGND.n407 117.001
R1084 VGND.n635 VGND.n479 117.001
R1085 VGND.n635 VGND.n473 117.001
R1086 VGND.n685 VGND.n684 117.001
R1087 VGND.n684 VGND.n454 117.001
R1088 VGND.n462 VGND.n461 117.001
R1089 VGND.n465 VGND.n462 117.001
R1090 VGND.n459 VGND.n458 117.001
R1091 VGND.n458 VGND.n450 117.001
R1092 VGND.n642 VGND.n641 117.001
R1093 VGND.n641 VGND.n450 117.001
R1094 VGND.n646 VGND.n645 117.001
R1095 VGND.n645 VGND.n454 117.001
R1096 VGND.n638 VGND.n637 117.001
R1097 VGND.n637 VGND.n473 117.001
R1098 VGND.n481 VGND.n480 117.001
R1099 VGND.n609 VGND.n481 117.001
R1100 VGND.n433 VGND.n413 117.001
R1101 VGND.n433 VGND.n407 117.001
R1102 VGND.n745 VGND.n744 117.001
R1103 VGND.n744 VGND.n284 117.001
R1104 VGND.n294 VGND.n293 117.001
R1105 VGND.n397 VGND.n294 117.001
R1106 VGND.n702 VGND.n701 117.001
R1107 VGND.n702 VGND.n281 117.001
R1108 VGND.n706 VGND.n705 117.001
R1109 VGND.n705 VGND.n281 117.001
R1110 VGND.n709 VGND.n292 117.001
R1111 VGND.n292 VGND.n284 117.001
R1112 VGND.n436 VGND.n435 117.001
R1113 VGND.n435 VGND.n407 117.001
R1114 VGND.n415 VGND.n414 117.001
R1115 VGND.n416 VGND.n415 117.001
R1116 VGND.n95 VGND.n94 117.001
R1117 VGND.n94 VGND.n66 117.001
R1118 VGND.n33 VGND.n31 117.001
R1119 VGND.n37 VGND.n33 117.001
R1120 VGND.n109 VGND.n108 117.001
R1121 VGND.n108 VGND.n37 117.001
R1122 VGND.n102 VGND.n96 117.001
R1123 VGND.n102 VGND.n34 117.001
R1124 VGND.n106 VGND.n105 117.001
R1125 VGND.n105 VGND.n34 117.001
R1126 VGND.n991 VGND.n55 117.001
R1127 VGND.n55 VGND.n53 117.001
R1128 VGND.n89 VGND.n87 117.001
R1129 VGND.n87 VGND.n78 117.001
R1130 VGND.n92 VGND.n91 117.001
R1131 VGND.n91 VGND.n66 117.001
R1132 VGND.n75 VGND.n74 117.001
R1133 VGND.n74 VGND.n66 117.001
R1134 VGND.n999 VGND.n998 117.001
R1135 VGND.n998 VGND.n37 117.001
R1136 VGND.n50 VGND.n46 117.001
R1137 VGND.n53 VGND.n46 117.001
R1138 VGND.n64 VGND.n60 117.001
R1139 VGND.n64 VGND.n34 117.001
R1140 VGND.n67 VGND.n61 117.001
R1141 VGND.n67 VGND.n34 117.001
R1142 VGND.n48 VGND.n45 117.001
R1143 VGND.n45 VGND.n37 117.001
R1144 VGND.n82 VGND.n81 117.001
R1145 VGND.n81 VGND.n66 117.001
R1146 VGND.n77 VGND.n76 117.001
R1147 VGND.n78 VGND.n77 117.001
R1148 VGND.n185 VGND.n184 117.001
R1149 VGND.n185 VGND.n180 117.001
R1150 VGND.n174 VGND.n136 117.001
R1151 VGND.n174 VGND.n11 117.001
R1152 VGND.n146 VGND.n138 117.001
R1153 VGND.n170 VGND.n138 117.001
R1154 VGND.n164 VGND 117.001
R1155 VGND.n164 VGND.n163 117.001
R1156 VGND.n157 VGND.n156 117.001
R1157 VGND.n156 VGND.n155 117.001
R1158 VGND VGND.n150 117.001
R1159 VGND.n162 VGND.n144 117.001
R1160 VGND.n163 VGND.n162 117.001
R1161 VGND.n169 VGND 117.001
R1162 VGND.n170 VGND.n169 117.001
R1163 VGND.n137 VGND 117.001
R1164 VGND.n137 VGND.n11 117.001
R1165 VGND.n238 VGND.n135 117.001
R1166 VGND.n179 VGND 117.001
R1167 VGND.n238 VGND.n179 117.001
R1168 VGND.n204 VGND.n203 117.001
R1169 VGND.n203 VGND.n187 117.001
R1170 VGND.n199 VGND.n190 117.001
R1171 VGND.n199 VGND.n187 117.001
R1172 VGND.n192 VGND.n191 117.001
R1173 VGND.n191 VGND.n181 117.001
R1174 VGND.n231 VGND.n182 117.001
R1175 VGND.n182 VGND.n181 117.001
R1176 VGND.n215 VGND.n214 117.001
R1177 VGND.n214 VGND.n196 117.001
R1178 VGND.n219 VGND.n218 117.001
R1179 VGND.n219 VGND.n196 117.001
R1180 VGND.n8 VGND.n6 117.001
R1181 VGND.n9 VGND.n8 117.001
R1182 VGND.n959 VGND.n956 117.001
R1183 VGND.n956 VGND.n17 117.001
R1184 VGND.n957 VGND.n955 117.001
R1185 VGND.n955 VGND.n17 117.001
R1186 VGND.n22 VGND.n20 117.001
R1187 VGND.n20 VGND.n17 117.001
R1188 VGND.n21 VGND.n19 117.001
R1189 VGND.n19 VGND.n17 117.001
R1190 VGND.n598 VGND.n587 117.001
R1191 VGND.n605 VGND.n587 117.001
R1192 VGND.n595 VGND.n593 117.001
R1193 VGND.n595 VGND.n260 117.001
R1194 VGND.n976 VGND.n975 117.001
R1195 VGND.n975 VGND.n974 117.001
R1196 VGND.n967 VGND.n966 117.001
R1197 VGND.n968 VGND.n967 117.001
R1198 VGND.n604 VGND.n603 117.001
R1199 VGND.n605 VGND.n604 117.001
R1200 VGND.n592 VGND.n591 117.001
R1201 VGND.n591 VGND.n260 117.001
R1202 VGND.n973 VGND.n972 117.001
R1203 VGND.n974 VGND.n973 117.001
R1204 VGND.n970 VGND.n969 117.001
R1205 VGND.n969 VGND.n968 117.001
R1206 VGND VGND.n760 115.576
R1207 VGND.n154 VGND.n150 109.642
R1208 VGND.n609 VGND.n608 108.163
R1209 VGND.n397 VGND.n396 108.163
R1210 VGND.n78 VGND.n16 108.163
R1211 VGND.n1024 VGND.n10 96.1003
R1212 VGND.n178 VGND.n177 93.2369
R1213 VGND.n235 VGND.n234 90.9521
R1214 VGND.n550 VGND.n502 90.3534
R1215 VGND.n555 VGND.n502 90.3534
R1216 VGND.n549 VGND.n512 90.3534
R1217 VGND.n544 VGND.n512 90.3534
R1218 VGND.n934 VGND.n776 90.3534
R1219 VGND.n776 VGND.n763 90.3534
R1220 VGND.n774 VGND.n773 90.3534
R1221 VGND.n773 VGND.n762 90.3534
R1222 VGND.n926 VGND.n830 90.3534
R1223 VGND.n834 VGND.n830 90.3534
R1224 VGND.n928 VGND.n829 90.3534
R1225 VGND.n832 VGND.n829 90.3534
R1226 VGND.n855 VGND.n854 90.3534
R1227 VGND.n854 VGND.n845 90.3534
R1228 VGND.n907 VGND.n844 90.3534
R1229 VGND.n912 VGND.n844 90.3534
R1230 VGND.n929 VGND.n826 89.9911
R1231 VGND VGND.n151 89.224
R1232 VGND VGND.n147 89.224
R1233 VGND.n158 VGND 89.224
R1234 VGND.n158 VGND.n157 89.224
R1235 VGND VGND.n143 89.224
R1236 VGND VGND.n168 89.224
R1237 VGND.n168 VGND.n144 89.224
R1238 VGND.n151 VGND.n144 89.224
R1239 VGND.n145 VGND.n136 89.224
R1240 VGND.n146 VGND.n145 89.224
R1241 VGND.n147 VGND.n146 89.224
R1242 VGND.n143 VGND 89.224
R1243 VGND.n734 VGND.n402 85.0829
R1244 VGND.n736 VGND.n401 85.0829
R1245 VGND.n719 VGND.n403 85.0829
R1246 VGND.n714 VGND.n425 85.0829
R1247 VGND.n425 VGND.n277 85.0829
R1248 VGND.n701 VGND.n289 85.0829
R1249 VGND.n706 VGND.n700 85.0829
R1250 VGND.n707 VGND.n706 85.0829
R1251 VGND.n728 VGND.n413 85.0829
R1252 VGND.n746 VGND.n745 85.0829
R1253 VGND.n460 VGND.n459 85.0829
R1254 VGND.n642 VGND.n446 85.0829
R1255 VGND.n643 VGND.n642 85.0829
R1256 VGND.n669 VGND.n479 85.0829
R1257 VGND.n686 VGND.n685 85.0829
R1258 VGND.n627 VGND.n625 85.0829
R1259 VGND.n660 VGND.n625 85.0829
R1260 VGND.n675 VGND.n469 85.0829
R1261 VGND.n677 VGND.n468 85.0829
R1262 VGND.n619 VGND.n470 85.0829
R1263 VGND.n201 VGND.n190 85.0829
R1264 VGND.n224 VGND.n192 85.0829
R1265 VGND.n192 VGND.n5 85.0829
R1266 VGND.n205 VGND.n204 85.0829
R1267 VGND.n216 VGND.n215 85.0829
R1268 VGND.n60 VGND.n42 85.0829
R1269 VGND.n127 VGND.n61 85.0829
R1270 VGND.n79 VGND.n61 85.0829
R1271 VGND.n121 VGND.n75 85.0829
R1272 VGND.n1000 VGND.n999 85.0829
R1273 VGND.n96 VGND.n30 85.0829
R1274 VGND.n112 VGND.n96 85.0829
R1275 VGND.n106 VGND.n101 85.0829
R1276 VGND.n109 VGND.n56 85.0829
R1277 VGND.n98 VGND.n95 85.0829
R1278 VGND.n116 VGND.n89 84.9588
R1279 VGND.n664 VGND.n615 84.9588
R1280 VGND.n723 VGND.n422 84.9588
R1281 VGND.n437 VGND.n414 84.9588
R1282 VGND.n633 VGND.n480 84.9588
R1283 VGND.n229 VGND.n184 84.9588
R1284 VGND.n84 VGND.n76 84.9588
R1285 VGND.n293 VGND.n272 84.6953
R1286 VGND.n737 VGND.n273 84.6953
R1287 VGND.n461 VGND.n441 84.6953
R1288 VGND.n678 VGND.n442 84.6953
R1289 VGND.n218 VGND.n2 84.6953
R1290 VGND.n51 VGND.n50 84.6953
R1291 VGND.n991 VGND.n990 84.6953
R1292 VGND.n964 VGND.n17 83.7263
R1293 VGND.n1020 VGND.n17 83.7263
R1294 VGND VGND.n929 77.2563
R1295 VGND.n720 VGND.n277 66.6518
R1296 VGND.n700 VGND.n698 66.6518
R1297 VGND.n631 VGND.n446 66.6518
R1298 VGND.n661 VGND.n660 66.6518
R1299 VGND.n225 VGND.n224 66.6518
R1300 VGND.n127 VGND.n126 66.6518
R1301 VGND.n113 VGND.n112 66.6518
R1302 VGND.n699 VGND.n291 64.7759
R1303 VGND.n751 VGND.n278 64.7759
R1304 VGND.n691 VGND.n447 64.7759
R1305 VGND.n659 VGND.n658 64.7759
R1306 VGND.n223 VGND.n194 64.7759
R1307 VGND.n128 VGND.n44 64.7759
R1308 VGND.n111 VGND.n110 64.7759
R1309 VGND.n700 VGND.n699 63.1207
R1310 VGND.n751 VGND.n277 63.1207
R1311 VGND.n691 VGND.n446 63.1207
R1312 VGND.n660 VGND.n659 63.1207
R1313 VGND.n224 VGND.n223 63.1207
R1314 VGND.n128 VGND.n127 63.1207
R1315 VGND.n112 VGND.n111 63.1207
R1316 VGND.n721 VGND.n720 61.2449
R1317 VGND.n698 VGND.n439 61.2449
R1318 VGND.n632 VGND.n631 61.2449
R1319 VGND.n662 VGND.n661 61.2449
R1320 VGND.n225 VGND.n183 61.2449
R1321 VGND.n126 VGND.n62 61.2449
R1322 VGND.n114 VGND.n113 61.2449
R1323 VGND.n549 VGND.n548 59.4829
R1324 VGND.n551 VGND.n549 59.4829
R1325 VGND.n551 VGND.n550 59.4829
R1326 VGND.n550 VGND.n501 59.4829
R1327 VGND.n920 VGND.n774 59.4829
R1328 VGND.n935 VGND.n774 59.4829
R1329 VGND.n935 VGND.n934 59.4829
R1330 VGND.n934 VGND.n933 59.4829
R1331 VGND.n835 VGND.n834 59.4829
R1332 VGND.n834 VGND.n833 59.4829
R1333 VGND.n833 VGND.n832 59.4829
R1334 VGND.n832 VGND.n831 59.4829
R1335 VGND.n894 VGND.n845 59.4829
R1336 VGND.n911 VGND.n845 59.4829
R1337 VGND.n912 VGND.n911 59.4829
R1338 VGND.n913 VGND.n912 59.4829
R1339 VGND.n401 VGND.n278 58.5793
R1340 VGND.n721 VGND.n719 58.5793
R1341 VGND.n439 VGND.n413 58.5793
R1342 VGND.n745 VGND.n291 58.5793
R1343 VGND.n632 VGND.n479 58.5793
R1344 VGND.n685 VGND.n447 58.5793
R1345 VGND.n658 VGND.n468 58.5793
R1346 VGND.n662 VGND.n619 58.5793
R1347 VGND.n204 VGND.n183 58.5793
R1348 VGND.n215 VGND.n194 58.5793
R1349 VGND.n75 VGND.n62 58.5793
R1350 VGND.n999 VGND.n44 58.5793
R1351 VGND.n110 VGND.n109 58.5793
R1352 VGND.n114 VGND.n95 58.5793
R1353 VGND.n402 VGND.n277 54.2123
R1354 VGND.n701 VGND.n700 54.2123
R1355 VGND.n459 VGND.n446 54.2123
R1356 VGND.n660 VGND.n469 54.2123
R1357 VGND.n224 VGND.n190 54.2123
R1358 VGND.n127 VGND.n60 54.2123
R1359 VGND.n112 VGND.n106 54.2123
R1360 VGND.n1023 VGND.n12 48.1018
R1361 VGND.n464 VGND.n442 41.7862
R1362 VGND.n681 VGND.n464 41.7862
R1363 VGND.n680 VGND.n679 41.7862
R1364 VGND.n681 VGND.n680 41.7862
R1365 VGND.n614 VGND.n611 41.7862
R1366 VGND.n666 VGND.n611 41.7862
R1367 VGND.n665 VGND.n664 41.7862
R1368 VGND.n666 VGND.n665 41.7862
R1369 VGND.n295 VGND.n273 41.7862
R1370 VGND.n741 VGND.n295 41.7862
R1371 VGND.n739 VGND.n738 41.7862
R1372 VGND.n741 VGND.n739 41.7862
R1373 VGND.n421 VGND.n418 41.7862
R1374 VGND.n725 VGND.n418 41.7862
R1375 VGND.n724 VGND.n723 41.7862
R1376 VGND.n725 VGND.n724 41.7862
R1377 VGND.n463 VGND.n441 41.7862
R1378 VGND.n681 VGND.n463 41.7862
R1379 VGND.n633 VGND.n610 41.7862
R1380 VGND.n666 VGND.n610 41.7862
R1381 VGND.n668 VGND.n667 41.7862
R1382 VGND.n667 VGND.n666 41.7862
R1383 VGND.n683 VGND.n682 41.7862
R1384 VGND.n682 VGND.n681 41.7862
R1385 VGND.n742 VGND.n272 41.7862
R1386 VGND.n742 VGND.n741 41.7862
R1387 VGND.n437 VGND.n417 41.7862
R1388 VGND.n725 VGND.n417 41.7862
R1389 VGND.n727 VGND.n726 41.7862
R1390 VGND.n726 VGND.n725 41.7862
R1391 VGND.n740 VGND.n290 41.7862
R1392 VGND.n741 VGND.n740 41.7862
R1393 VGND.n990 VGND.n52 41.7862
R1394 VGND.n995 VGND.n52 41.7862
R1395 VGND.n993 VGND.n992 41.7862
R1396 VGND.n995 VGND.n993 41.7862
R1397 VGND.n97 VGND.n86 41.7862
R1398 VGND.n118 VGND.n86 41.7862
R1399 VGND.n117 VGND.n116 41.7862
R1400 VGND.n118 VGND.n117 41.7862
R1401 VGND.n996 VGND.n51 41.7862
R1402 VGND.n996 VGND.n995 41.7862
R1403 VGND.n85 VGND.n84 41.7862
R1404 VGND.n118 VGND.n85 41.7862
R1405 VGND.n120 VGND.n119 41.7862
R1406 VGND.n119 VGND.n118 41.7862
R1407 VGND.n994 VGND.n43 41.7862
R1408 VGND.n995 VGND.n994 41.7862
R1409 VGND.n229 VGND.n228 41.7862
R1410 VGND.n228 VGND.n227 41.7862
R1411 VGND.n207 VGND.n206 41.7862
R1412 VGND.n208 VGND.n207 41.7862
R1413 VGND.n220 VGND.n2 41.7862
R1414 VGND.n221 VGND.n220 41.7862
R1415 VGND.n217 VGND.n197 41.7862
R1416 VGND.n211 VGND.n197 41.7862
R1417 VGND VGND.n544 40.4485
R1418 VGND.n555 VGND 40.4485
R1419 VGND VGND.n555 40.4485
R1420 VGND VGND.n762 40.4485
R1421 VGND VGND.n763 40.4485
R1422 VGND VGND.n763 40.4485
R1423 VGND VGND.n855 40.4485
R1424 VGND VGND.n907 40.4485
R1425 VGND.n907 VGND 40.4485
R1426 VGND.n544 VGND.n503 38.1445
R1427 VGND.n939 VGND.n762 38.1445
R1428 VGND.n906 VGND.n855 38.1445
R1429 VGND.n661 VGND.n476 34.4123
R1430 VGND.n672 VGND.n476 34.4123
R1431 VGND.n659 VGND.n453 34.4123
R1432 VGND.n689 VGND.n453 34.4123
R1433 VGND.n676 VGND.n455 34.4123
R1434 VGND.n689 VGND.n455 34.4123
R1435 VGND.n674 VGND.n673 34.4123
R1436 VGND.n673 VGND.n672 34.4123
R1437 VGND.n626 VGND.n475 34.4123
R1438 VGND.n672 VGND.n475 34.4123
R1439 VGND.n652 VGND.n452 34.4123
R1440 VGND.n689 VGND.n452 34.4123
R1441 VGND.n720 VGND.n410 34.4123
R1442 VGND.n731 VGND.n410 34.4123
R1443 VGND.n751 VGND.n750 34.4123
R1444 VGND.n750 VGND.n749 34.4123
R1445 VGND.n735 VGND.n285 34.4123
R1446 VGND.n749 VGND.n285 34.4123
R1447 VGND.n733 VGND.n732 34.4123
R1448 VGND.n732 VGND.n731 34.4123
R1449 VGND.n715 VGND.n409 34.4123
R1450 VGND.n731 VGND.n409 34.4123
R1451 VGND.n429 VGND.n283 34.4123
R1452 VGND.n749 VGND.n283 34.4123
R1453 VGND.n631 VGND.n477 34.4123
R1454 VGND.n672 VGND.n477 34.4123
R1455 VGND.n691 VGND.n690 34.4123
R1456 VGND.n690 VGND.n689 34.4123
R1457 VGND.n647 VGND.n451 34.4123
R1458 VGND.n689 VGND.n451 34.4123
R1459 VGND.n639 VGND.n474 34.4123
R1460 VGND.n672 VGND.n474 34.4123
R1461 VGND.n671 VGND.n670 34.4123
R1462 VGND.n672 VGND.n671 34.4123
R1463 VGND.n688 VGND.n687 34.4123
R1464 VGND.n689 VGND.n688 34.4123
R1465 VGND.n698 VGND.n411 34.4123
R1466 VGND.n731 VGND.n411 34.4123
R1467 VGND.n699 VGND.n286 34.4123
R1468 VGND.n749 VGND.n286 34.4123
R1469 VGND.n710 VGND.n282 34.4123
R1470 VGND.n749 VGND.n282 34.4123
R1471 VGND.n432 VGND.n408 34.4123
R1472 VGND.n731 VGND.n408 34.4123
R1473 VGND.n730 VGND.n729 34.4123
R1474 VGND.n731 VGND.n730 34.4123
R1475 VGND.n748 VGND.n747 34.4123
R1476 VGND.n749 VGND.n748 34.4123
R1477 VGND.n113 VGND.n71 34.4123
R1478 VGND.n124 VGND.n71 34.4123
R1479 VGND.n111 VGND.n36 34.4123
R1480 VGND.n1003 VGND.n36 34.4123
R1481 VGND.n100 VGND.n38 34.4123
R1482 VGND.n1003 VGND.n38 34.4123
R1483 VGND.n99 VGND.n72 34.4123
R1484 VGND.n124 VGND.n72 34.4123
R1485 VGND.n90 VGND.n70 34.4123
R1486 VGND.n124 VGND.n70 34.4123
R1487 VGND.n1005 VGND.n1004 34.4123
R1488 VGND.n1004 VGND.n1003 34.4123
R1489 VGND.n126 VGND.n125 34.4123
R1490 VGND.n125 VGND.n124 34.4123
R1491 VGND.n128 VGND.n39 34.4123
R1492 VGND.n1003 VGND.n39 34.4123
R1493 VGND.n47 VGND.n35 34.4123
R1494 VGND.n1003 VGND.n35 34.4123
R1495 VGND.n80 VGND.n69 34.4123
R1496 VGND.n124 VGND.n69 34.4123
R1497 VGND.n123 VGND.n122 34.4123
R1498 VGND.n124 VGND.n123 34.4123
R1499 VGND.n1002 VGND.n1001 34.4123
R1500 VGND.n1003 VGND.n1002 34.4123
R1501 VGND.n241 VGND.n240 34.4123
R1502 VGND.n240 VGND.n239 34.4123
R1503 VGND.n236 VGND.n134 34.4123
R1504 VGND.n237 VGND.n236 34.4123
R1505 VGND.n226 VGND.n225 34.4123
R1506 VGND.n227 VGND.n226 34.4123
R1507 VGND.n233 VGND.n232 34.4123
R1508 VGND.n234 VGND.n233 34.4123
R1509 VGND.n209 VGND.n202 34.4123
R1510 VGND.n209 VGND.n208 34.4123
R1511 VGND.n223 VGND.n222 34.4123
R1512 VGND.n222 VGND.n221 34.4123
R1513 VGND.n1027 VGND.n1026 34.4123
R1514 VGND.n1026 VGND.n1025 34.4123
R1515 VGND.n212 VGND.n198 34.4123
R1516 VGND.n212 VGND.n211 34.4123
R1517 VGND.n352 VGND.n347 32.5005
R1518 VGND.n353 VGND.n352 32.5005
R1519 VGND.n357 VGND 32.5005
R1520 VGND.n357 VGND.n12 32.5005
R1521 VGND.n354 VGND 32.5005
R1522 VGND.n354 VGND.n353 32.5005
R1523 VGND.n363 VGND.n362 32.5005
R1524 VGND.n363 VGND.n12 32.5005
R1525 VGND.n367 VGND 32.5005
R1526 VGND.n367 VGND.n366 32.5005
R1527 VGND.n373 VGND.n372 32.5005
R1528 VGND.n374 VGND.n373 32.5005
R1529 VGND.n365 VGND.n340 32.5005
R1530 VGND.n366 VGND.n365 32.5005
R1531 VGND VGND.n332 32.5005
R1532 VGND.n374 VGND.n332 32.5005
R1533 VGND.n338 VGND.n337 32.5005
R1534 VGND.n337 VGND.n325 32.5005
R1535 VGND VGND.n324 32.5005
R1536 VGND.n383 VGND.n324 32.5005
R1537 VGND VGND.n378 32.5005
R1538 VGND.n378 VGND.n325 32.5005
R1539 VGND.n384 VGND.n323 32.5005
R1540 VGND.n384 VGND.n383 32.5005
R1541 VGND.n388 VGND 32.5005
R1542 VGND.n388 VGND.n387 32.5005
R1543 VGND.n394 VGND.n393 32.5005
R1544 VGND.n395 VGND.n394 32.5005
R1545 VGND.n386 VGND.n302 32.5005
R1546 VGND.n387 VGND.n386 32.5005
R1547 VGND VGND.n297 32.5005
R1548 VGND.n395 VGND.n297 32.5005
R1549 VGND.n314 VGND.n313 32.5005
R1550 VGND.n315 VGND.n314 32.5005
R1551 VGND VGND.n268 32.5005
R1552 VGND.n268 VGND.n266 32.5005
R1553 VGND VGND.n316 32.5005
R1554 VGND.n316 VGND.n315 32.5005
R1555 VGND.n269 VGND.n267 32.5005
R1556 VGND.n267 VGND.n266 32.5005
R1557 VGND.n350 VGND.n349 19.5005
R1558 VGND.n351 VGND.n349 19.5005
R1559 VGND.n360 VGND.n359 19.5005
R1560 VGND.n359 VGND.n13 19.5005
R1561 VGND.n355 VGND.n344 19.5005
R1562 VGND.n344 VGND.n343 19.5005
R1563 VGND.n370 VGND.n369 19.5005
R1564 VGND.n369 VGND.n335 19.5005
R1565 VGND.n376 VGND.n334 19.5005
R1566 VGND.n376 VGND.n375 19.5005
R1567 VGND.n381 VGND.n380 19.5005
R1568 VGND.n382 VGND.n381 19.5005
R1569 VGND.n329 VGND.n321 19.5005
R1570 VGND.n321 VGND.n320 19.5005
R1571 VGND.n391 VGND.n390 19.5005
R1572 VGND.n390 VGND.n298 19.5005
R1573 VGND.n306 VGND.n303 19.5005
R1574 VGND.n306 VGND.n296 19.5005
R1575 VGND.n311 VGND.n310 19.5005
R1576 VGND.n310 VGND.n308 19.5005
R1577 VGND.n950 VGND.n949 19.5005
R1578 VGND.n951 VGND.n950 19.5005
R1579 VGND.n426 VGND.n278 18.297
R1580 VGND.n722 VGND.n721 18.297
R1581 VGND.n439 VGND.n438 18.297
R1582 VGND.n708 VGND.n291 18.297
R1583 VGND.n634 VGND.n632 18.297
R1584 VGND.n644 VGND.n447 18.297
R1585 VGND.n658 VGND.n657 18.297
R1586 VGND.n663 VGND.n662 18.297
R1587 VGND.n230 VGND.n183 18.297
R1588 VGND.n194 VGND.n193 18.297
R1589 VGND.n83 VGND.n62 18.297
R1590 VGND.n49 VGND.n44 18.297
R1591 VGND.n110 VGND.n57 18.297
R1592 VGND.n115 VGND.n114 18.297
R1593 VGND.n172 VGND.n140 17.2064
R1594 VGND.n172 VGND.n171 17.2064
R1595 VGND.n167 VGND.n166 17.2064
R1596 VGND.n166 VGND.n141 17.2064
R1597 VGND.n160 VGND.n159 17.2064
R1598 VGND.n160 VGND.n149 17.2064
R1599 VGND.n153 VGND.n152 17.2064
R1600 VGND.n176 VGND.n175 17.2064
R1601 VGND.n175 VGND.n10 17.2064
R1602 VGND.n116 VGND.n115 8.08353
R1603 VGND.n664 VGND.n663 8.08353
R1604 VGND.n723 VGND.n722 8.08353
R1605 VGND.n426 VGND.n273 8.08353
R1606 VGND.n438 VGND.n437 8.08353
R1607 VGND.n708 VGND.n272 8.08353
R1608 VGND.n634 VGND.n633 8.08353
R1609 VGND.n644 VGND.n441 8.08353
R1610 VGND.n657 VGND.n442 8.08353
R1611 VGND.n230 VGND.n229 8.08353
R1612 VGND.n193 VGND.n2 8.08353
R1613 VGND.n84 VGND.n83 8.08353
R1614 VGND.n51 VGND.n49 8.08353
R1615 VGND.n990 VGND.n57 8.08353
R1616 VGND.n1014 VGND.n1013 6.64112
R1617 VGND.n155 VGND.n154 5.84938
R1618 VGND.n535 VGND.n495 5.57862
R1619 VGND.n942 VGND.n759 5.57706
R1620 VGND.n533 VGND 5.02361
R1621 VGND.n761 VGND 5.02361
R1622 VGND.n761 VGND 5.02361
R1623 VGND.n904 VGND 5.02361
R1624 VGND.n532 VGND 5.01717
R1625 VGND.n537 VGND 5.01717
R1626 VGND.n494 VGND 5.01717
R1627 VGND.n494 VGND 5.01717
R1628 VGND.n580 VGND 5.01717
R1629 VGND.n580 VGND 5.01717
R1630 VGND.n870 VGND 5.01717
R1631 VGND.n870 VGND 5.01717
R1632 VGND.n903 VGND 5.01717
R1633 VGND.n903 VGND 5.01717
R1634 VGND.n797 VGND 5.01717
R1635 VGND.n797 VGND 5.01717
R1636 VGND.n807 VGND 5.01717
R1637 VGND.n807 VGND 5.01717
R1638 VGND.n1015 VGND 5.01717
R1639 VGND.n1016 VGND 5.01717
R1640 VGND.n254 VGND 5.01717
R1641 VGND.n254 VGND 5.01717
R1642 VGND.n600 VGND 5.01717
R1643 VGND.n600 VGND 5.01717
R1644 VGND.n757 VGND 5.00093
R1645 VGND.n247 VGND 4.25376
R1646 VGND.n250 VGND 3.49683
R1647 VGND.n1037 VGND 3.37909
R1648 VGND.n752 VGND.n276 3.27485
R1649 VGND.n692 VGND.n445 3.27485
R1650 VGND.n129 VGND.n26 3.27485
R1651 VGND.n58 VGND.n27 3.27485
R1652 VGND.n620 VGND.n443 3.27485
R1653 VGND.n697 VGND.n274 3.27485
R1654 VGND.n189 VGND.n3 3.27485
R1655 VGND.n428 VGND.n426 3.08756
R1656 VGND.n722 VGND.n717 3.08756
R1657 VGND.n438 VGND.n436 3.08756
R1658 VGND.n709 VGND.n708 3.08756
R1659 VGND.n638 VGND.n634 3.08756
R1660 VGND.n646 VGND.n644 3.08756
R1661 VGND.n657 VGND.n656 3.08756
R1662 VGND.n663 VGND.n617 3.08756
R1663 VGND.n231 VGND.n230 3.08756
R1664 VGND.n193 VGND.n6 3.08756
R1665 VGND.n83 VGND.n82 3.08756
R1666 VGND.n49 VGND.n48 3.08756
R1667 VGND.n57 VGND.n31 3.08756
R1668 VGND.n115 VGND.n92 3.08756
R1669 VGND.n440 VGND 3.06629
R1670 VGND.n629 VGND 3.06629
R1671 VGND.n1009 VGND 3.06629
R1672 VGND.n927 VGND 3.01226
R1673 VGND.n270 VGND 2.51601
R1674 VGND.n980 VGND.n979 2.46929
R1675 VGND.n949 VGND.n948 2.35839
R1676 VGND VGND.n503 2.3045
R1677 VGND.n939 VGND 2.3045
R1678 VGND VGND.n906 2.3045
R1679 VGND.n270 VGND 2.11902
R1680 VGND.n1013 VGND.n24 1.98151
R1681 VGND.n532 VGND.n531 1.96988
R1682 VGND.n431 VGND 1.91991
R1683 VGND.n649 VGND 1.91991
R1684 VGND.n29 VGND 1.91991
R1685 VGND.n581 VGND.n579 1.8605
R1686 VGND.n539 VGND.n538 1.8605
R1687 VGND.n568 VGND.n567 1.8605
R1688 VGND.n582 VGND.n581 1.8605
R1689 VGND.n567 VGND.n566 1.8605
R1690 VGND.n902 VGND.n856 1.8605
R1691 VGND.n818 VGND.n817 1.8605
R1692 VGND.n808 VGND.n806 1.8605
R1693 VGND.n879 VGND.n878 1.8605
R1694 VGND.n902 VGND.n901 1.8605
R1695 VGND.n819 VGND.n818 1.8605
R1696 VGND.n809 VGND.n808 1.8605
R1697 VGND.n878 VGND.n877 1.8605
R1698 VGND.n958 VGND.n23 1.8605
R1699 VGND.n1018 VGND.n1017 1.8605
R1700 VGND.n978 VGND.n255 1.8605
R1701 VGND.n601 VGND.n599 1.8605
R1702 VGND.n978 VGND.n977 1.8605
R1703 VGND.n602 VGND.n601 1.8605
R1704 VGND.n943 VGND.n942 1.79344
R1705 VGND.n535 VGND.n249 1.68993
R1706 VGND.n130 VGND.n58 1.55665
R1707 VGND.n693 VGND.n443 1.55665
R1708 VGND.n753 VGND.n274 1.55665
R1709 VGND.n753 VGND.n752 1.55665
R1710 VGND.n693 VGND.n692 1.55665
R1711 VGND.n1032 VGND.n3 1.55665
R1712 VGND.n130 VGND.n129 1.55665
R1713 VGND.n1010 VGND.n27 1.43327
R1714 VGND.n628 VGND.n620 1.43327
R1715 VGND.n697 VGND.n696 1.43327
R1716 VGND.n696 VGND.n276 1.43327
R1717 VGND.n628 VGND.n445 1.43327
R1718 VGND.n189 VGND.n133 1.43327
R1719 VGND.n1010 VGND.n26 1.43327
R1720 VGND.n243 VGND.n134 1.21955
R1721 VGND.n130 VGND 0.946224
R1722 VGND.n693 VGND 0.946224
R1723 VGND.n753 VGND 0.946224
R1724 VGND.n430 VGND 0.905763
R1725 VGND.n630 VGND 0.905763
R1726 VGND.n1008 VGND 0.905763
R1727 VGND.n754 VGND.n272 0.846996
R1728 VGND.n754 VGND.n273 0.846996
R1729 VGND.n694 VGND.n441 0.846996
R1730 VGND.n694 VGND.n442 0.846996
R1731 VGND.n1033 VGND.n2 0.846996
R1732 VGND.n989 VGND.n51 0.846996
R1733 VGND.n990 VGND.n989 0.846996
R1734 VGND VGND.n536 0.827844
R1735 VGND VGND 0.771099
R1736 VGND.n1012 VGND.n25 0.760382
R1737 VGND.n534 VGND.n503 0.715885
R1738 VGND.n906 VGND.n905 0.715885
R1739 VGND.n940 VGND.n760 0.715885
R1740 VGND.n940 VGND.n939 0.715885
R1741 VGND.n1030 VGND 0.695143
R1742 VGND.n699 VGND.n274 0.664786
R1743 VGND.n698 VGND.n697 0.664786
R1744 VGND.n752 VGND.n751 0.664786
R1745 VGND.n720 VGND.n276 0.664786
R1746 VGND.n692 VGND.n691 0.664786
R1747 VGND.n631 VGND.n445 0.664786
R1748 VGND.n659 VGND.n443 0.664786
R1749 VGND.n661 VGND.n620 0.664786
R1750 VGND.n223 VGND.n3 0.664786
R1751 VGND.n225 VGND.n189 0.664786
R1752 VGND.n245 VGND 0.664786
R1753 VGND.n129 VGND.n128 0.664786
R1754 VGND.n126 VGND.n26 0.664786
R1755 VGND.n111 VGND.n58 0.664786
R1756 VGND.n113 VGND.n27 0.664786
R1757 VGND.n4 VGND 0.644695
R1758 VGND.n758 VGND.n247 0.64299
R1759 VGND VGND 0.635531
R1760 VGND.n250 VGND.n248 0.629595
R1761 VGND.n241 VGND.n177 0.582318
R1762 VGND.n253 VGND.n24 0.568833
R1763 VGND.n252 VGND.n25 0.568833
R1764 VGND.n244 VGND.n243 0.517167
R1765 VGND VGND 0.457722
R1766 VGND.n59 VGND 0.447211
R1767 VGND.n444 VGND 0.447211
R1768 VGND.n275 VGND 0.447211
R1769 VGND.n696 VGND 0.439349
R1770 VGND.n628 VGND 0.439349
R1771 VGND.n1010 VGND 0.439349
R1772 VGND VGND 0.406319
R1773 VGND.n905 VGND 0.405187
R1774 VGND.n941 VGND.n940 0.402844
R1775 VGND.n536 VGND.n534 0.401281
R1776 VGND.n695 VGND.n246 0.393625
R1777 VGND.n987 VGND.n986 0.393625
R1778 VGND.n602 VGND 0.376971
R1779 VGND.n977 VGND 0.376971
R1780 VGND.n599 VGND 0.376971
R1781 VGND.n582 VGND 0.376971
R1782 VGND.n568 VGND 0.376971
R1783 VGND.n539 VGND 0.376971
R1784 VGND.n531 VGND 0.376971
R1785 VGND.n579 VGND 0.376971
R1786 VGND.n566 VGND 0.376971
R1787 VGND VGND.n809 0.376971
R1788 VGND VGND.n819 0.376971
R1789 VGND.n901 VGND 0.376971
R1790 VGND.n879 VGND 0.376971
R1791 VGND.n806 VGND 0.376971
R1792 VGND.n817 VGND 0.376971
R1793 VGND VGND.n856 0.376971
R1794 VGND.n927 VGND.n760 0.376971
R1795 VGND.n877 VGND 0.376971
R1796 VGND.n714 VGND.n713 0.376971
R1797 VGND.n711 VGND.n707 0.376971
R1798 VGND.n648 VGND.n643 0.376971
R1799 VGND.n651 VGND.n627 0.376971
R1800 VGND.n1028 VGND.n5 0.376971
R1801 VGND.n79 VGND.n28 0.376971
R1802 VGND VGND.n1018 0.376971
R1803 VGND.n958 VGND 0.376971
R1804 VGND.n1006 VGND.n30 0.376971
R1805 VGND VGND.n255 0.376971
R1806 VGND.n534 VGND.n533 0.376281
R1807 VGND.n905 VGND.n904 0.376281
R1808 VGND.n940 VGND.n761 0.376281
R1809 VGND.n252 VGND.n251 0.365484
R1810 VGND.n1011 VGND.n1010 0.346566
R1811 VGND.n1032 VGND 0.342762
R1812 VGND.n59 VGND.n29 0.321553
R1813 VGND.n649 VGND.n444 0.321553
R1814 VGND.n431 VGND.n275 0.321553
R1815 VGND.n440 VGND.n430 0.321553
R1816 VGND.n630 VGND.n629 0.321553
R1817 VGND.n1009 VGND.n1008 0.321553
R1818 VGND.n1031 VGND 0.318384
R1819 VGND.n948 VGND.n947 0.304262
R1820 VGND.n986 VGND.n985 0.285503
R1821 VGND.n757 VGND.n246 0.279901
R1822 VGND.n943 VGND.n249 0.250766
R1823 VGND.n980 VGND.n253 0.247336
R1824 VGND.n944 VGND 0.233324
R1825 VGND.n1031 VGND.n1030 0.228964
R1826 VGND.n947 VGND.n271 0.218382
R1827 VGND.n986 VGND.n0 0.209183
R1828 VGND.n1017 VGND 0.208833
R1829 VGND.n946 VGND 0.203416
R1830 VGND.n1035 VGND.n1 0.203021
R1831 VGND.n981 VGND.n249 0.200936
R1832 VGND.n985 VGND.n246 0.196464
R1833 VGND.n271 VGND.n270 0.188289
R1834 VGND.n712 VGND.n430 0.186355
R1835 VGND.n650 VGND.n630 0.186355
R1836 VGND.n1008 VGND.n1007 0.186355
R1837 VGND.n756 VGND.n755 0.181262
R1838 VGND.n1035 VGND.n1034 0.181262
R1839 VGND.n130 VGND.n59 0.171553
R1840 VGND.n693 VGND.n444 0.171553
R1841 VGND.n753 VGND.n275 0.171553
R1842 VGND.n947 VGND.n946 0.169234
R1843 VGND.n988 VGND 0.166889
R1844 VGND.n567 VGND 0.166125
R1845 VGND.n818 VGND 0.166125
R1846 VGND.n538 VGND 0.164562
R1847 VGND.n581 VGND 0.164562
R1848 VGND.n902 VGND 0.164562
R1849 VGND.n808 VGND 0.164562
R1850 VGND.n601 VGND 0.164562
R1851 VGND.n712 VGND.n431 0.158395
R1852 VGND.n650 VGND.n649 0.158395
R1853 VGND.n1007 VGND.n29 0.158395
R1854 VGND.n1011 VGND.n23 0.14931
R1855 VGND.n696 VGND.n440 0.145237
R1856 VGND.n629 VGND.n628 0.145237
R1857 VGND.n1010 VGND.n1009 0.145237
R1858 VGND.n1036 VGND.n1035 0.144712
R1859 VGND.n1017 VGND.n1016 0.139389
R1860 VGND.n756 VGND.n1 0.137606
R1861 VGND.n713 VGND.n712 0.133357
R1862 VGND.n712 VGND.n711 0.133357
R1863 VGND.n650 VGND.n648 0.133357
R1864 VGND.n651 VGND.n650 0.133357
R1865 VGND.n1029 VGND.n1028 0.133357
R1866 VGND.n1007 VGND.n28 0.133357
R1867 VGND.n1007 VGND.n1006 0.133357
R1868 VGND VGND.n4 0.126904
R1869 VGND.n982 VGND.n981 0.126796
R1870 VGND.n695 VGND 0.124938
R1871 VGND VGND.n988 0.123766
R1872 VGND.n271 VGND 0.111032
R1873 VGND.n1014 VGND.n23 0.110619
R1874 VGND.n538 VGND.n537 0.109875
R1875 VGND.n581 VGND.n580 0.109875
R1876 VGND.n878 VGND.n870 0.109875
R1877 VGND.n903 VGND.n902 0.109875
R1878 VGND.n808 VGND.n807 0.109875
R1879 VGND.n601 VGND.n600 0.109875
R1880 VGND.n132 VGND 0.10256
R1881 VGND.n758 VGND 0.0991948
R1882 VGND.n567 VGND.n495 0.0934687
R1883 VGND.n1012 VGND.n1011 0.0907506
R1884 VGND.n818 VGND.n759 0.0903438
R1885 VGND.n979 VGND.n254 0.0860255
R1886 VGND.n248 VGND 0.0836655
R1887 VGND.n1033 VGND.n1032 0.0803611
R1888 VGND.n536 VGND.n535 0.0780862
R1889 VGND.n942 VGND.n941 0.0780862
R1890 VGND.n1013 VGND.n1012 0.0780862
R1891 VGND.n133 VGND 0.0759438
R1892 VGND VGND.n1015 0.0699444
R1893 VGND.n1016 VGND 0.0699444
R1894 VGND.n985 VGND.n984 0.0687
R1895 VGND VGND.n1037 0.0686031
R1896 VGND.n1029 VGND.n4 0.0677619
R1897 VGND.n754 VGND.n753 0.0651358
R1898 VGND.n694 VGND.n693 0.0651358
R1899 VGND VGND.n694 0.0651358
R1900 VGND.n989 VGND.n130 0.0651358
R1901 VGND.n989 VGND 0.0651358
R1902 VGND.n1032 VGND.n1031 0.0624048
R1903 VGND.n1034 VGND 0.0620278
R1904 VGND.n1030 VGND.n1029 0.0576429
R1905 VGND.n755 VGND 0.0572671
R1906 VGND VGND.n532 0.0551875
R1907 VGND.n537 VGND 0.0551875
R1908 VGND.n494 VGND 0.0551875
R1909 VGND.n580 VGND 0.0551875
R1910 VGND.n870 VGND 0.0551875
R1911 VGND VGND.n903 0.0551875
R1912 VGND VGND.n797 0.0551875
R1913 VGND.n807 VGND 0.0551875
R1914 VGND VGND.n254 0.0551875
R1915 VGND.n600 VGND 0.0551875
R1916 VGND.n131 VGND 0.0524663
R1917 VGND.n981 VGND.n980 0.0501588
R1918 VGND.n983 VGND.n1 0.0478611
R1919 VGND.n533 VGND 0.0434688
R1920 VGND.n904 VGND 0.0434688
R1921 VGND VGND.n761 0.0434688
R1922 VGND.n131 VGND 0.0433241
R1923 VGND.n696 VGND.n695 0.042429
R1924 VGND.n132 VGND.n131 0.0417809
R1925 VGND.n133 VGND.n132 0.0416985
R1926 VGND VGND 0.0346797
R1927 VGND.n987 VGND.n245 0.0316884
R1928 VGND.n1011 VGND 0.0297969
R1929 VGND.n988 VGND.n987 0.0294694
R1930 VGND.n1015 VGND.n1014 0.0292698
R1931 VGND.n979 VGND.n978 0.0233551
R1932 VGND.n797 VGND.n759 0.0200312
R1933 VGND.n1034 VGND.n1033 0.0188333
R1934 VGND.n495 VGND.n494 0.0169062
R1935 VGND.n946 VGND.n945 0.0134167
R1936 VGND.n244 VGND.n133 0.0120878
R1937 VGND.n253 VGND.n252 0.010792
R1938 VGND VGND.n756 0.00952437
R1939 VGND.n755 VGND.n754 0.00836871
R1940 VGND VGND.n943 0.00513139
R1941 VGND.n25 VGND.n24 0.00492478
R1942 VGND.n941 VGND 0.00284375
R1943 VGND.n984 VGND.n247 0.00178858
R1944 VGND.n982 VGND.n248 0.00173884
R1945 VGND.n1037 VGND.n1036 0.00165108
R1946 VGND.n251 VGND.n250 0.00164397
R1947 VGND.n944 VGND.n758 0.00129115
R1948 VGND.n245 VGND.n244 0.000993097
R1949 VGND.n945 VGND.n944 0.00073924
R1950 VGND.n251 VGND.n0 0.000549738
R1951 VGND.n983 VGND.n982 0.000530793
R1952 VGND.n1036 VGND.n0 0.000528422
R1953 VGND.n984 VGND.n983 0.00051895
R1954 VGND.n945 VGND.n757 0.000514212
R1955 VDPWR.n451 VDPWR.n340 5809.41
R1956 VDPWR.n340 VDPWR.n336 5809.41
R1957 VDPWR.n424 VDPWR.n360 5809.41
R1958 VDPWR.n424 VDPWR.n361 5809.41
R1959 VDPWR.n286 VDPWR.n138 5809.41
R1960 VDPWR.n286 VDPWR.n139 5809.41
R1961 VDPWR.n244 VDPWR.n145 5809.41
R1962 VDPWR.n163 VDPWR.n145 5809.41
R1963 VDPWR.n289 VDPWR.n288 5809.41
R1964 VDPWR.n288 VDPWR.n134 5809.41
R1965 VDPWR.n255 VDPWR.n146 5809.41
R1966 VDPWR.n255 VDPWR.n147 5809.41
R1967 VDPWR.n630 VDPWR.n581 5809.41
R1968 VDPWR.n631 VDPWR.n630 5809.41
R1969 VDPWR.n430 VDPWR.n429 5784.71
R1970 VDPWR.n429 VDPWR.n358 5784.71
R1971 VDPWR.n368 VDPWR.n365 5784.71
R1972 VDPWR.n419 VDPWR.n365 5784.71
R1973 VDPWR.n273 VDPWR.n268 5784.71
R1974 VDPWR.n269 VDPWR.n268 5784.71
R1975 VDPWR.n248 VDPWR.n157 5784.71
R1976 VDPWR.n157 VDPWR.n155 5784.71
R1977 VDPWR.n266 VDPWR.n257 5784.71
R1978 VDPWR.n266 VDPWR.n258 5784.71
R1979 VDPWR.n154 VDPWR.n151 5784.71
R1980 VDPWR.n250 VDPWR.n151 5784.71
R1981 VDPWR.n595 VDPWR.n592 5784.71
R1982 VDPWR.n595 VDPWR.n580 5784.71
R1983 VDPWR.n388 VDPWR.n384 4912.94
R1984 VDPWR.n400 VDPWR.n384 4912.94
R1985 VDPWR.n388 VDPWR.n385 4912.94
R1986 VDPWR.n400 VDPWR.n385 4912.94
R1987 VDPWR.n344 VDPWR.n343 4912.94
R1988 VDPWR.n448 VDPWR.n343 4912.94
R1989 VDPWR.n447 VDPWR.n344 4912.94
R1990 VDPWR.n448 VDPWR.n447 4912.94
R1991 VDPWR.n168 VDPWR.n165 4912.94
R1992 VDPWR.n241 VDPWR.n165 4912.94
R1993 VDPWR.n168 VDPWR.n166 4912.94
R1994 VDPWR.n241 VDPWR.n166 4912.94
R1995 VDPWR.n303 VDPWR.n120 4912.94
R1996 VDPWR.n282 VDPWR.n120 4912.94
R1997 VDPWR.n303 VDPWR.n121 4912.94
R1998 VDPWR.n282 VDPWR.n121 4912.94
R1999 VDPWR.n215 VDPWR.n193 4912.94
R2000 VDPWR.n215 VDPWR.n164 4912.94
R2001 VDPWR.n206 VDPWR.n193 4912.94
R2002 VDPWR.n206 VDPWR.n164 4912.94
R2003 VDPWR.n301 VDPWR.n123 4912.94
R2004 VDPWR.n280 VDPWR.n123 4912.94
R2005 VDPWR.n301 VDPWR.n124 4912.94
R2006 VDPWR.n280 VDPWR.n124 4912.94
R2007 VDPWR.n585 VDPWR.n584 4912.94
R2008 VDPWR.n609 VDPWR.n584 4912.94
R2009 VDPWR.n606 VDPWR.n585 4912.94
R2010 VDPWR.n609 VDPWR.n606 4912.94
R2011 VDPWR.n627 VDPWR.n613 4912.94
R2012 VDPWR.n618 VDPWR.n614 4912.94
R2013 VDPWR.n627 VDPWR.n614 4912.94
R2014 VDPWR.n444 VDPWR.n348 4207.06
R2015 VDPWR.n348 VDPWR.n347 4207.06
R2016 VDPWR.n454 VDPWR.n333 4207.06
R2017 VDPWR.n335 VDPWR.n333 4207.06
R2018 VDPWR.n416 VDPWR.n372 4207.06
R2019 VDPWR.n372 VDPWR.n369 4207.06
R2020 VDPWR.n404 VDPWR.n377 4207.06
R2021 VDPWR.n383 VDPWR.n377 4207.06
R2022 VDPWR.n307 VDPWR.n111 4207.06
R2023 VDPWR.n309 VDPWR.n111 4207.06
R2024 VDPWR.n315 VDPWR.n107 4207.06
R2025 VDPWR.n107 VDPWR.n103 4207.06
R2026 VDPWR.n203 VDPWR.n202 4207.06
R2027 VDPWR.n202 VDPWR.n195 4207.06
R2028 VDPWR.n221 VDPWR.n220 4207.06
R2029 VDPWR.n222 VDPWR.n221 4207.06
R2030 VDPWR.n126 VDPWR.n116 4207.06
R2031 VDPWR.n126 VDPWR.n114 4207.06
R2032 VDPWR.n317 VDPWR.n101 4207.06
R2033 VDPWR.n104 VDPWR.n101 4207.06
R2034 VDPWR.n179 VDPWR.n171 4207.06
R2035 VDPWR.n232 VDPWR.n171 4207.06
R2036 VDPWR.n229 VDPWR.n173 4207.06
R2037 VDPWR.n230 VDPWR.n229 4207.06
R2038 VDPWR.n603 VDPWR.n589 4207.06
R2039 VDPWR.n589 VDPWR.n588 4207.06
R2040 VDPWR.n638 VDPWR.n569 4207.06
R2041 VDPWR.n640 VDPWR.n569 4207.06
R2042 VDPWR.n430 VDPWR.n338 4020
R2043 VDPWR.n358 VDPWR.n350 4020
R2044 VDPWR.n378 VDPWR.n368 4020
R2045 VDPWR.n419 VDPWR.n366 4020
R2046 VDPWR.n273 VDPWR.n272 4020
R2047 VDPWR.n270 VDPWR.n269 4020
R2048 VDPWR.n248 VDPWR.n158 4020
R2049 VDPWR.n211 VDPWR.n155 4020
R2050 VDPWR.n257 VDPWR.n133 4020
R2051 VDPWR.n260 VDPWR.n258 4020
R2052 VDPWR.n207 VDPWR.n154 4020
R2053 VDPWR.n250 VDPWR.n152 4020
R2054 VDPWR.n592 VDPWR.n579 4020
R2055 VDPWR.n632 VDPWR.n580 4020
R2056 VDPWR.n451 VDPWR.n338 3998.82
R2057 VDPWR.n350 VDPWR.n336 3998.82
R2058 VDPWR.n378 VDPWR.n360 3998.82
R2059 VDPWR.n366 VDPWR.n361 3998.82
R2060 VDPWR.n272 VDPWR.n138 3998.82
R2061 VDPWR.n270 VDPWR.n139 3998.82
R2062 VDPWR.n244 VDPWR.n158 3998.82
R2063 VDPWR.n211 VDPWR.n163 3998.82
R2064 VDPWR.n289 VDPWR.n133 3998.82
R2065 VDPWR.n260 VDPWR.n134 3998.82
R2066 VDPWR.n207 VDPWR.n146 3998.82
R2067 VDPWR.n152 VDPWR.n147 3998.82
R2068 VDPWR.n581 VDPWR.n579 3998.82
R2069 VDPWR.n632 VDPWR.n631 3998.82
R2070 VDPWR.n444 VDPWR.n332 3409.41
R2071 VDPWR.n454 VDPWR.n332 3409.41
R2072 VDPWR.n433 VDPWR.n347 3409.41
R2073 VDPWR.n433 VDPWR.n335 3409.41
R2074 VDPWR.n416 VDPWR.n373 3409.41
R2075 VDPWR.n404 VDPWR.n373 3409.41
R2076 VDPWR.n382 VDPWR.n369 3409.41
R2077 VDPWR.n383 VDPWR.n382 3409.41
R2078 VDPWR.n307 VDPWR.n106 3409.41
R2079 VDPWR.n315 VDPWR.n106 3409.41
R2080 VDPWR.n310 VDPWR.n309 3409.41
R2081 VDPWR.n310 VDPWR.n103 3409.41
R2082 VDPWR.n203 VDPWR.n187 3409.41
R2083 VDPWR.n220 VDPWR.n187 3409.41
R2084 VDPWR.n195 VDPWR.n186 3409.41
R2085 VDPWR.n222 VDPWR.n186 3409.41
R2086 VDPWR.n116 VDPWR.n100 3409.41
R2087 VDPWR.n317 VDPWR.n100 3409.41
R2088 VDPWR.n293 VDPWR.n114 3409.41
R2089 VDPWR.n293 VDPWR.n104 3409.41
R2090 VDPWR.n179 VDPWR.n178 3409.41
R2091 VDPWR.n178 VDPWR.n173 3409.41
R2092 VDPWR.n232 VDPWR.n231 3409.41
R2093 VDPWR.n231 VDPWR.n230 3409.41
R2094 VDPWR.n603 VDPWR.n572 3409.41
R2095 VDPWR.n638 VDPWR.n572 3409.41
R2096 VDPWR.n588 VDPWR.n568 3409.41
R2097 VDPWR.n640 VDPWR.n568 3409.41
R2098 VDPWR.n698 VDPWR.n683 1789.41
R2099 VDPWR.n705 VDPWR.n683 1789.41
R2100 VDPWR.n698 VDPWR.n684 1789.41
R2101 VDPWR.n705 VDPWR.n684 1789.41
R2102 VDPWR.n714 VDPWR.n676 1789.41
R2103 VDPWR.n695 VDPWR.n676 1789.41
R2104 VDPWR.n714 VDPWR.n677 1789.41
R2105 VDPWR.n695 VDPWR.n677 1789.41
R2106 VDPWR.n826 VDPWR.n819 1789.41
R2107 VDPWR.n819 VDPWR.n817 1789.41
R2108 VDPWR.n838 VDPWR.n671 1789.41
R2109 VDPWR.n840 VDPWR.n671 1789.41
R2110 VDPWR.n800 VDPWR.n781 1789.41
R2111 VDPWR.n800 VDPWR.n782 1789.41
R2112 VDPWR.n814 VDPWR.n740 1789.41
R2113 VDPWR.n814 VDPWR.n741 1789.41
R2114 VDPWR.n774 VDPWR.n746 1789.41
R2115 VDPWR.n803 VDPWR.n746 1789.41
R2116 VDPWR.n774 VDPWR.n747 1789.41
R2117 VDPWR.n803 VDPWR.n747 1789.41
R2118 VDPWR.n766 VDPWR.n758 1789.41
R2119 VDPWR.n758 VDPWR.n753 1789.41
R2120 VDPWR.n766 VDPWR.n759 1789.41
R2121 VDPWR.n759 VDPWR.n753 1789.41
R2122 VDPWR.n700 VDPWR.n686 1789.41
R2123 VDPWR.n703 VDPWR.n686 1789.41
R2124 VDPWR.n700 VDPWR.n687 1789.41
R2125 VDPWR.n703 VDPWR.n687 1789.41
R2126 VDPWR.n689 VDPWR.n674 1789.41
R2127 VDPWR.n694 VDPWR.n689 1789.41
R2128 VDPWR.n690 VDPWR.n674 1789.41
R2129 VDPWR.n694 VDPWR.n690 1789.41
R2130 VDPWR.n818 VDPWR.n737 1789.41
R2131 VDPWR.n828 VDPWR.n737 1789.41
R2132 VDPWR.n733 VDPWR.n717 1789.41
R2133 VDPWR.n733 VDPWR.n673 1789.41
R2134 VDPWR.n776 VDPWR.n749 1789.41
R2135 VDPWR.n779 VDPWR.n749 1789.41
R2136 VDPWR.n776 VDPWR.n750 1789.41
R2137 VDPWR.n779 VDPWR.n750 1789.41
R2138 VDPWR.n768 VDPWR.n754 1789.41
R2139 VDPWR.n771 VDPWR.n754 1789.41
R2140 VDPWR.n768 VDPWR.n755 1789.41
R2141 VDPWR.n771 VDPWR.n755 1789.41
R2142 VDPWR.n505 VDPWR.n479 1789.41
R2143 VDPWR.n479 VDPWR.n475 1789.41
R2144 VDPWR.n505 VDPWR.n480 1789.41
R2145 VDPWR.n480 VDPWR.n475 1789.41
R2146 VDPWR.n478 VDPWR.n472 1789.41
R2147 VDPWR.n507 VDPWR.n472 1789.41
R2148 VDPWR.n478 VDPWR.n473 1789.41
R2149 VDPWR.n507 VDPWR.n473 1789.41
R2150 VDPWR.n488 VDPWR.n483 1789.41
R2151 VDPWR.n497 VDPWR.n483 1789.41
R2152 VDPWR.n488 VDPWR.n484 1789.41
R2153 VDPWR.n497 VDPWR.n484 1789.41
R2154 VDPWR.n490 VDPWR.n486 1789.41
R2155 VDPWR.n495 VDPWR.n490 1789.41
R2156 VDPWR.n491 VDPWR.n486 1789.41
R2157 VDPWR.n495 VDPWR.n491 1789.41
R2158 VDPWR.n553 VDPWR.n527 1789.41
R2159 VDPWR.n527 VDPWR.n523 1789.41
R2160 VDPWR.n553 VDPWR.n528 1789.41
R2161 VDPWR.n528 VDPWR.n523 1789.41
R2162 VDPWR.n526 VDPWR.n520 1789.41
R2163 VDPWR.n555 VDPWR.n520 1789.41
R2164 VDPWR.n526 VDPWR.n521 1789.41
R2165 VDPWR.n555 VDPWR.n521 1789.41
R2166 VDPWR.n536 VDPWR.n531 1789.41
R2167 VDPWR.n545 VDPWR.n531 1789.41
R2168 VDPWR.n536 VDPWR.n532 1789.41
R2169 VDPWR.n545 VDPWR.n532 1789.41
R2170 VDPWR.n538 VDPWR.n534 1789.41
R2171 VDPWR.n543 VDPWR.n538 1789.41
R2172 VDPWR.n539 VDPWR.n534 1789.41
R2173 VDPWR.n543 VDPWR.n539 1789.41
R2174 VDPWR.n354 VDPWR.n338 1789.41
R2175 VDPWR.n354 VDPWR.n350 1789.41
R2176 VDPWR.n379 VDPWR.n378 1789.41
R2177 VDPWR.n379 VDPWR.n366 1789.41
R2178 VDPWR.n82 VDPWR.n5 1789.41
R2179 VDPWR.n85 VDPWR.n5 1789.41
R2180 VDPWR.n83 VDPWR.n82 1789.41
R2181 VDPWR.n76 VDPWR.n9 1789.41
R2182 VDPWR.n79 VDPWR.n9 1789.41
R2183 VDPWR.n76 VDPWR.n10 1789.41
R2184 VDPWR.n79 VDPWR.n10 1789.41
R2185 VDPWR.n56 VDPWR.n27 1789.41
R2186 VDPWR.n54 VDPWR.n27 1789.41
R2187 VDPWR.n73 VDPWR.n14 1789.41
R2188 VDPWR.n73 VDPWR.n15 1789.41
R2189 VDPWR.n48 VDPWR.n29 1789.41
R2190 VDPWR.n51 VDPWR.n29 1789.41
R2191 VDPWR.n48 VDPWR.n30 1789.41
R2192 VDPWR.n51 VDPWR.n30 1789.41
R2193 VDPWR.n45 VDPWR.n34 1789.41
R2194 VDPWR.n42 VDPWR.n35 1789.41
R2195 VDPWR.n45 VDPWR.n35 1789.41
R2196 VDPWR.n272 VDPWR.n271 1789.41
R2197 VDPWR.n271 VDPWR.n270 1789.41
R2198 VDPWR.n212 VDPWR.n158 1789.41
R2199 VDPWR.n212 VDPWR.n211 1789.41
R2200 VDPWR.n261 VDPWR.n133 1789.41
R2201 VDPWR.n261 VDPWR.n260 1789.41
R2202 VDPWR.n208 VDPWR.n207 1789.41
R2203 VDPWR.n208 VDPWR.n152 1789.41
R2204 VDPWR.n633 VDPWR.n579 1789.41
R2205 VDPWR.n633 VDPWR.n632 1789.41
R2206 VDPWR.n628 VDPWR.n612 1534.21
R2207 VDPWR VDPWR.n616 1446.4
R2208 VDPWR.n619 VDPWR 1446.4
R2209 VDPWR.n53 VDPWR.n52 1315.04
R2210 VDPWR.n719 VDPWR.n718 1231.76
R2211 VDPWR.n718 VDPWR.n670 1231.76
R2212 VDPWR.n821 VDPWR.n721 1231.76
R2213 VDPWR.n821 VDPWR.n820 1231.76
R2214 VDPWR.n790 VDPWR.n789 1231.76
R2215 VDPWR.n789 VDPWR.n788 1231.76
R2216 VDPWR.n795 VDPWR.n784 1231.76
R2217 VDPWR.n795 VDPWR.n785 1231.76
R2218 VDPWR.n729 VDPWR.n726 1231.76
R2219 VDPWR.n729 VDPWR.n728 1231.76
R2220 VDPWR.n830 VDPWR.n725 1231.76
R2221 VDPWR.n830 VDPWR.n829 1231.76
R2222 VDPWR.n25 VDPWR.n24 1231.76
R2223 VDPWR.n24 VDPWR.n20 1231.76
R2224 VDPWR.n58 VDPWR.n23 1231.76
R2225 VDPWR.n58 VDPWR.n19 1231.76
R2226 VDPWR.n618 VDPWR.n617 1189.42
R2227 VDPWR.n434 VDPWR.n332 797.648
R2228 VDPWR.n434 VDPWR.n433 797.648
R2229 VDPWR.n381 VDPWR.n373 797.648
R2230 VDPWR.n382 VDPWR.n381 797.648
R2231 VDPWR.n311 VDPWR.n106 797.648
R2232 VDPWR.n311 VDPWR.n310 797.648
R2233 VDPWR.n210 VDPWR.n187 797.648
R2234 VDPWR.n210 VDPWR.n186 797.648
R2235 VDPWR.n294 VDPWR.n100 797.648
R2236 VDPWR.n294 VDPWR.n293 797.648
R2237 VDPWR.n178 VDPWR.n172 797.648
R2238 VDPWR.n231 VDPWR.n172 797.648
R2239 VDPWR.n573 VDPWR.n572 797.648
R2240 VDPWR.n573 VDPWR.n568 797.648
R2241 VDPWR.n826 VDPWR.n721 557.648
R2242 VDPWR.n836 VDPWR.n721 557.648
R2243 VDPWR.n836 VDPWR.n719 557.648
R2244 VDPWR.n838 VDPWR.n719 557.648
R2245 VDPWR.n820 VDPWR.n817 557.648
R2246 VDPWR.n820 VDPWR.n723 557.648
R2247 VDPWR.n723 VDPWR.n670 557.648
R2248 VDPWR.n840 VDPWR.n670 557.648
R2249 VDPWR.n784 VDPWR.n781 557.648
R2250 VDPWR.n792 VDPWR.n784 557.648
R2251 VDPWR.n792 VDPWR.n790 557.648
R2252 VDPWR.n790 VDPWR.n740 557.648
R2253 VDPWR.n785 VDPWR.n782 557.648
R2254 VDPWR.n786 VDPWR.n785 557.648
R2255 VDPWR.n788 VDPWR.n786 557.648
R2256 VDPWR.n788 VDPWR.n741 557.648
R2257 VDPWR.n818 VDPWR.n725 557.648
R2258 VDPWR.n834 VDPWR.n725 557.648
R2259 VDPWR.n834 VDPWR.n726 557.648
R2260 VDPWR.n726 VDPWR.n717 557.648
R2261 VDPWR.n829 VDPWR.n828 557.648
R2262 VDPWR.n829 VDPWR.n724 557.648
R2263 VDPWR.n728 VDPWR.n724 557.648
R2264 VDPWR.n728 VDPWR.n673 557.648
R2265 VDPWR.n56 VDPWR.n23 557.648
R2266 VDPWR.n68 VDPWR.n23 557.648
R2267 VDPWR.n68 VDPWR.n25 557.648
R2268 VDPWR.n25 VDPWR.n14 557.648
R2269 VDPWR.n54 VDPWR.n19 557.648
R2270 VDPWR.n70 VDPWR.n19 557.648
R2271 VDPWR.n70 VDPWR.n20 557.648
R2272 VDPWR.n20 VDPWR.n15 557.648
R2273 VDPWR.n626 VDPWR.n615 524.069
R2274 VDPWR.n629 VDPWR.n628 473.772
R2275 VDPWR.n626 VDPWR.n625 473.219
R2276 VDPWR.n352 VDPWR.n351 447.06
R2277 VDPWR.n423 VDPWR.n422 447.06
R2278 VDPWR.n245 VDPWR.n161 447.06
R2279 VDPWR.n285 VDPWR.n276 447.06
R2280 VDPWR.n259 VDPWR.n136 447.06
R2281 VDPWR.n254 VDPWR.n253 447.06
R2282 VDPWR.n583 VDPWR.n582 447.06
R2283 VDPWR.n357 VDPWR.n349 444.515
R2284 VDPWR.n420 VDPWR.n364 444.515
R2285 VDPWR.n247 VDPWR.n159 444.515
R2286 VDPWR.n274 VDPWR.n143 444.515
R2287 VDPWR.n265 VDPWR.n264 444.515
R2288 VDPWR.n251 VDPWR.n150 444.515
R2289 VDPWR.n596 VDPWR.n591 444.515
R2290 VDPWR.n616 VDPWR.n615 432.942
R2291 VDPWR.n357 VDPWR.n356 428.8
R2292 VDPWR.n421 VDPWR.n420 428.8
R2293 VDPWR.n247 VDPWR.n246 428.8
R2294 VDPWR.n275 VDPWR.n274 428.8
R2295 VDPWR.n264 VDPWR.n263 428.8
R2296 VDPWR.n252 VDPWR.n251 428.8
R2297 VDPWR.n591 VDPWR.n578 428.8
R2298 VDPWR.n356 VDPWR.n352 426.541
R2299 VDPWR.n422 VDPWR.n421 426.541
R2300 VDPWR.n246 VDPWR.n245 426.541
R2301 VDPWR.n276 VDPWR.n275 426.541
R2302 VDPWR.n263 VDPWR.n259 426.541
R2303 VDPWR.n253 VDPWR.n252 426.541
R2304 VDPWR.n582 VDPWR.n578 426.541
R2305 VDPWR.n620 VDPWR.n619 387.368
R2306 VDPWR.n443 VDPWR.n330 363.671
R2307 VDPWR.n415 VDPWR.n414 363.671
R2308 VDPWR.n198 VDPWR.n184 363.671
R2309 VDPWR.n112 VDPWR.n110 363.671
R2310 VDPWR.n125 VDPWR.n98 363.671
R2311 VDPWR.n181 VDPWR.n180 363.671
R2312 VDPWR.n597 VDPWR.n566 363.671
R2313 VDPWR.n456 VDPWR.n455 363.295
R2314 VDPWR.n413 VDPWR.n405 363.295
R2315 VDPWR.n224 VDPWR.n223 363.295
R2316 VDPWR.n277 VDPWR.n94 363.295
R2317 VDPWR.n319 VDPWR.n318 363.295
R2318 VDPWR.n227 VDPWR.n226 363.295
R2319 VDPWR.n642 VDPWR.n641 363.295
R2320 VDPWR.n415 VDPWR.n374 362.37
R2321 VDPWR.n443 VDPWR.n442 362.37
R2322 VDPWR.n199 VDPWR.n198 362.37
R2323 VDPWR.n180 VDPWR.n177 362.37
R2324 VDPWR.n118 VDPWR.n112 362.37
R2325 VDPWR.n127 VDPWR.n125 362.37
R2326 VDPWR.n598 VDPWR.n597 362.37
R2327 VDPWR.n405 VDPWR.n376 361.584
R2328 VDPWR.n455 VDPWR.n331 361.584
R2329 VDPWR.n223 VDPWR.n185 361.584
R2330 VDPWR.n228 VDPWR.n227 361.584
R2331 VDPWR.n278 VDPWR.n277 361.584
R2332 VDPWR.n318 VDPWR.n99 361.584
R2333 VDPWR.n641 VDPWR.n567 361.584
R2334 VDPWR.n403 VDPWR.n380 349.733
R2335 VDPWR.n453 VDPWR.n334 349.733
R2336 VDPWR.n639 VDPWR.n570 349.733
R2337 VDPWR.n417 VDPWR.n370 341.769
R2338 VDPWR.n446 VDPWR.n445 341.769
R2339 VDPWR.n605 VDPWR.n604 341.769
R2340 VDPWR.n428 VDPWR.n425 304.478
R2341 VDPWR.n401 VDPWR.n359 285.291
R2342 VDPWR.n339 VDPWR.n337 285.291
R2343 VDPWR.n611 VDPWR.n610 285.291
R2344 VDPWR.n371 VDPWR.n367 269.361
R2345 VDPWR.n427 VDPWR.n426 269.361
R2346 VDPWR.n594 VDPWR.n593 269.361
R2347 VDPWR.n697 VDPWR 190.871
R2348 VDPWR.n706 VDPWR 190.871
R2349 VDPWR.n697 VDPWR.n682 190.871
R2350 VDPWR.n713 VDPWR 190.871
R2351 VDPWR.n678 VDPWR 190.871
R2352 VDPWR.n713 VDPWR.n712 190.871
R2353 VDPWR VDPWR.n825 190.871
R2354 VDPWR.n825 VDPWR.n824 190.871
R2355 VDPWR VDPWR.n669 190.871
R2356 VDPWR.n841 VDPWR.n669 190.871
R2357 VDPWR.n799 VDPWR 190.871
R2358 VDPWR.n799 VDPWR.n798 190.871
R2359 VDPWR.n813 VDPWR 190.871
R2360 VDPWR.n813 VDPWR.n812 190.871
R2361 VDPWR.n773 VDPWR 190.871
R2362 VDPWR.n804 VDPWR 190.871
R2363 VDPWR.n773 VDPWR.n745 190.871
R2364 VDPWR.n765 VDPWR 190.871
R2365 VDPWR.n760 VDPWR 190.871
R2366 VDPWR.n765 VDPWR.n764 190.871
R2367 VDPWR.n701 VDPWR.n688 190.871
R2368 VDPWR VDPWR.n701 190.871
R2369 VDPWR.n702 VDPWR 190.871
R2370 VDPWR.n692 VDPWR.n691 190.871
R2371 VDPWR VDPWR.n692 190.871
R2372 VDPWR.n693 VDPWR 190.871
R2373 VDPWR.n738 VDPWR.n727 190.871
R2374 VDPWR VDPWR.n738 190.871
R2375 VDPWR.n734 VDPWR.n732 190.871
R2376 VDPWR VDPWR.n734 190.871
R2377 VDPWR.n777 VDPWR.n751 190.871
R2378 VDPWR VDPWR.n777 190.871
R2379 VDPWR.n778 VDPWR 190.871
R2380 VDPWR.n770 VDPWR 190.871
R2381 VDPWR VDPWR.n769 190.871
R2382 VDPWR.n769 VDPWR.n757 190.871
R2383 VDPWR.n504 VDPWR 190.871
R2384 VDPWR.n481 VDPWR 190.871
R2385 VDPWR.n504 VDPWR.n503 190.871
R2386 VDPWR.n477 VDPWR 190.871
R2387 VDPWR.n508 VDPWR 190.871
R2388 VDPWR.n477 VDPWR.n471 190.871
R2389 VDPWR.n487 VDPWR.n482 190.871
R2390 VDPWR.n487 VDPWR 190.871
R2391 VDPWR.n498 VDPWR 190.871
R2392 VDPWR.n494 VDPWR 190.871
R2393 VDPWR VDPWR.n493 190.871
R2394 VDPWR.n493 VDPWR.n492 190.871
R2395 VDPWR.n552 VDPWR 190.871
R2396 VDPWR.n529 VDPWR 190.871
R2397 VDPWR.n552 VDPWR.n551 190.871
R2398 VDPWR.n525 VDPWR 190.871
R2399 VDPWR.n556 VDPWR 190.871
R2400 VDPWR.n525 VDPWR.n519 190.871
R2401 VDPWR.n535 VDPWR.n530 190.871
R2402 VDPWR.n535 VDPWR 190.871
R2403 VDPWR.n546 VDPWR 190.871
R2404 VDPWR.n542 VDPWR 190.871
R2405 VDPWR VDPWR.n541 190.871
R2406 VDPWR.n541 VDPWR.n540 190.871
R2407 VDPWR.n355 VDPWR.n353 190.871
R2408 VDPWR.n356 VDPWR.n355 190.871
R2409 VDPWR.n396 VDPWR.n363 190.871
R2410 VDPWR.n421 VDPWR.n363 190.871
R2411 VDPWR.n7 VDPWR.n4 190.871
R2412 VDPWR.n7 VDPWR 190.871
R2413 VDPWR.n86 VDPWR 190.871
R2414 VDPWR.n77 VDPWR.n12 190.871
R2415 VDPWR VDPWR.n77 190.871
R2416 VDPWR.n78 VDPWR 190.871
R2417 VDPWR.n57 VDPWR.n26 190.871
R2418 VDPWR VDPWR.n26 190.871
R2419 VDPWR.n72 VDPWR.n16 190.871
R2420 VDPWR.n72 VDPWR 190.871
R2421 VDPWR.n49 VDPWR.n32 190.871
R2422 VDPWR VDPWR.n49 190.871
R2423 VDPWR.n50 VDPWR 190.871
R2424 VDPWR.n44 VDPWR 190.871
R2425 VDPWR VDPWR.n43 190.871
R2426 VDPWR.n43 VDPWR.n40 190.871
R2427 VDPWR.n246 VDPWR.n160 190.871
R2428 VDPWR.n217 VDPWR.n160 190.871
R2429 VDPWR.n275 VDPWR.n142 190.871
R2430 VDPWR.n142 VDPWR.n141 190.871
R2431 VDPWR.n262 VDPWR.n131 190.871
R2432 VDPWR.n263 VDPWR.n262 190.871
R2433 VDPWR.n237 VDPWR.n149 190.871
R2434 VDPWR.n252 VDPWR.n149 190.871
R2435 VDPWR.n634 VDPWR.n578 190.871
R2436 VDPWR.n635 VDPWR.n634 190.871
R2437 VDPWR.n707 VDPWR.n706 190.494
R2438 VDPWR.n711 VDPWR.n678 190.494
R2439 VDPWR.n805 VDPWR.n804 190.494
R2440 VDPWR.n763 VDPWR.n760 190.494
R2441 VDPWR.n702 VDPWR.n680 190.494
R2442 VDPWR.n693 VDPWR.n679 190.494
R2443 VDPWR.n778 VDPWR.n744 190.494
R2444 VDPWR.n770 VDPWR.n756 190.494
R2445 VDPWR.n502 VDPWR.n481 190.494
R2446 VDPWR.n509 VDPWR.n508 190.494
R2447 VDPWR.n499 VDPWR.n498 190.494
R2448 VDPWR.n494 VDPWR.n469 190.494
R2449 VDPWR.n550 VDPWR.n529 190.494
R2450 VDPWR.n557 VDPWR.n556 190.494
R2451 VDPWR.n547 VDPWR.n546 190.494
R2452 VDPWR.n542 VDPWR.n517 190.494
R2453 VDPWR.n87 VDPWR.n86 190.494
R2454 VDPWR.n78 VDPWR.n11 190.494
R2455 VDPWR.n50 VDPWR.n31 190.494
R2456 VDPWR.n44 VDPWR.n39 190.494
R2457 VDPWR.n46 VDPWR.n33 179.118
R2458 VDPWR.n47 VDPWR.n28 179.118
R2459 VDPWR.n52 VDPWR.n28 179.118
R2460 VDPWR.n55 VDPWR.n53 179.118
R2461 VDPWR.n55 VDPWR.n21 179.118
R2462 VDPWR.n69 VDPWR.n21 179.118
R2463 VDPWR.n69 VDPWR.n22 179.118
R2464 VDPWR.n22 VDPWR.n13 179.118
R2465 VDPWR.n74 VDPWR.n13 179.118
R2466 VDPWR.n75 VDPWR.n8 179.118
R2467 VDPWR.n80 VDPWR.n8 179.118
R2468 VDPWR.n81 VDPWR.n6 179.118
R2469 VDPWR.n213 VDPWR.n162 174.868
R2470 VDPWR.n316 VDPWR.n102 174.868
R2471 VDPWR.n42 VDPWR.n41 173.642
R2472 VDPWR.n85 VDPWR.n84 173.642
R2473 VDPWR.n214 VDPWR.n156 170.885
R2474 VDPWR.n308 VDPWR.n115 170.885
R2475 VDPWR.n267 VDPWR.n256 152.239
R2476 VDPWR.n242 VDPWR.n144 142.645
R2477 VDPWR.n281 VDPWR.n137 142.645
R2478 VDPWR.n340 VDPWR.n339 137.326
R2479 VDPWR.n371 VDPWR.n365 136.964
R2480 VDPWR.n595 VDPWR.n594 136.964
R2481 VDPWR.n201 VDPWR.n153 134.68
R2482 VDPWR.n302 VDPWR.n122 134.68
R2483 VDPWR.n837 VDPWR.n668 131.388
R2484 VDPWR.n842 VDPWR.n668 131.388
R2485 VDPWR.n822 VDPWR.n720 131.388
R2486 VDPWR.n823 VDPWR.n822 131.388
R2487 VDPWR.n791 VDPWR.n742 131.388
R2488 VDPWR.n811 VDPWR.n742 131.388
R2489 VDPWR.n796 VDPWR.n783 131.388
R2490 VDPWR.n797 VDPWR.n796 131.388
R2491 VDPWR.n731 VDPWR.n730 131.388
R2492 VDPWR.n735 VDPWR.n730 131.388
R2493 VDPWR.n832 VDPWR.n831 131.388
R2494 VDPWR.n831 VDPWR.n736 131.388
R2495 VDPWR.n61 VDPWR.n17 131.388
R2496 VDPWR.n71 VDPWR.n17 131.388
R2497 VDPWR.n60 VDPWR.n59 131.388
R2498 VDPWR.n59 VDPWR.n18 131.388
R2499 VDPWR.n425 VDPWR.n359 123.096
R2500 VDPWR.n629 VDPWR.n611 123.096
R2501 VDPWR.n428 VDPWR.n427 122.733
R2502 VDPWR.n75 VDPWR.n74 120.168
R2503 VDPWR.n47 VDPWR.n46 117.9
R2504 VDPWR.n81 VDPWR.n80 117.9
R2505 VDPWR VDPWR.n616 97.577
R2506 VDPWR.n619 VDPWR 97.5373
R2507 VDPWR VDPWR.n750 92.5005
R2508 VDPWR.n750 VDPWR.n748 92.5005
R2509 VDPWR.n751 VDPWR.n749 92.5005
R2510 VDPWR.n749 VDPWR.n748 92.5005
R2511 VDPWR VDPWR.n673 92.5005
R2512 VDPWR.n839 VDPWR.n673 92.5005
R2513 VDPWR VDPWR.n724 92.5005
R2514 VDPWR.n835 VDPWR.n724 92.5005
R2515 VDPWR.n828 VDPWR 92.5005
R2516 VDPWR.n828 VDPWR.n827 92.5005
R2517 VDPWR.n818 VDPWR.n727 92.5005
R2518 VDPWR.n827 VDPWR.n818 92.5005
R2519 VDPWR.n834 VDPWR.n833 92.5005
R2520 VDPWR.n835 VDPWR.n834 92.5005
R2521 VDPWR.n732 VDPWR.n717 92.5005
R2522 VDPWR.n839 VDPWR.n717 92.5005
R2523 VDPWR VDPWR.n690 92.5005
R2524 VDPWR.n690 VDPWR.n675 92.5005
R2525 VDPWR.n691 VDPWR.n689 92.5005
R2526 VDPWR.n689 VDPWR.n675 92.5005
R2527 VDPWR VDPWR.n687 92.5005
R2528 VDPWR.n687 VDPWR.n685 92.5005
R2529 VDPWR.n688 VDPWR.n686 92.5005
R2530 VDPWR.n686 VDPWR.n685 92.5005
R2531 VDPWR.n764 VDPWR.n759 92.5005
R2532 VDPWR.n759 VDPWR.n752 92.5005
R2533 VDPWR VDPWR.n758 92.5005
R2534 VDPWR.n758 VDPWR.n752 92.5005
R2535 VDPWR.n747 VDPWR.n745 92.5005
R2536 VDPWR.n748 VDPWR.n747 92.5005
R2537 VDPWR.n746 VDPWR 92.5005
R2538 VDPWR.n748 VDPWR.n746 92.5005
R2539 VDPWR.n812 VDPWR.n741 92.5005
R2540 VDPWR.n741 VDPWR.n739 92.5005
R2541 VDPWR.n786 VDPWR.n743 92.5005
R2542 VDPWR.n793 VDPWR.n786 92.5005
R2543 VDPWR.n798 VDPWR.n782 92.5005
R2544 VDPWR.n782 VDPWR.n780 92.5005
R2545 VDPWR VDPWR.n781 92.5005
R2546 VDPWR.n781 VDPWR.n780 92.5005
R2547 VDPWR.n792 VDPWR 92.5005
R2548 VDPWR.n793 VDPWR.n792 92.5005
R2549 VDPWR VDPWR.n740 92.5005
R2550 VDPWR.n740 VDPWR.n739 92.5005
R2551 VDPWR.n841 VDPWR.n840 92.5005
R2552 VDPWR.n840 VDPWR.n839 92.5005
R2553 VDPWR.n723 VDPWR.n667 92.5005
R2554 VDPWR.n835 VDPWR.n723 92.5005
R2555 VDPWR.n824 VDPWR.n817 92.5005
R2556 VDPWR.n827 VDPWR.n817 92.5005
R2557 VDPWR.n826 VDPWR 92.5005
R2558 VDPWR.n827 VDPWR.n826 92.5005
R2559 VDPWR VDPWR.n836 92.5005
R2560 VDPWR.n836 VDPWR.n835 92.5005
R2561 VDPWR.n838 VDPWR 92.5005
R2562 VDPWR.n839 VDPWR.n838 92.5005
R2563 VDPWR.n712 VDPWR.n677 92.5005
R2564 VDPWR.n677 VDPWR.n675 92.5005
R2565 VDPWR VDPWR.n676 92.5005
R2566 VDPWR.n676 VDPWR.n675 92.5005
R2567 VDPWR.n684 VDPWR.n682 92.5005
R2568 VDPWR.n685 VDPWR.n684 92.5005
R2569 VDPWR.n683 VDPWR 92.5005
R2570 VDPWR.n685 VDPWR.n683 92.5005
R2571 VDPWR VDPWR.n755 92.5005
R2572 VDPWR.n755 VDPWR.n752 92.5005
R2573 VDPWR.n757 VDPWR.n754 92.5005
R2574 VDPWR.n754 VDPWR.n752 92.5005
R2575 VDPWR.n484 VDPWR 92.5005
R2576 VDPWR.n489 VDPWR.n484 92.5005
R2577 VDPWR.n483 VDPWR.n482 92.5005
R2578 VDPWR.n485 VDPWR.n483 92.5005
R2579 VDPWR.n473 VDPWR.n471 92.5005
R2580 VDPWR.n476 VDPWR.n473 92.5005
R2581 VDPWR.n472 VDPWR 92.5005
R2582 VDPWR.n474 VDPWR.n472 92.5005
R2583 VDPWR.n503 VDPWR.n480 92.5005
R2584 VDPWR.n480 VDPWR.n476 92.5005
R2585 VDPWR VDPWR.n479 92.5005
R2586 VDPWR.n479 VDPWR.n474 92.5005
R2587 VDPWR VDPWR.n491 92.5005
R2588 VDPWR.n491 VDPWR.n489 92.5005
R2589 VDPWR.n492 VDPWR.n490 92.5005
R2590 VDPWR.n490 VDPWR.n485 92.5005
R2591 VDPWR.n532 VDPWR 92.5005
R2592 VDPWR.n537 VDPWR.n532 92.5005
R2593 VDPWR.n531 VDPWR.n530 92.5005
R2594 VDPWR.n533 VDPWR.n531 92.5005
R2595 VDPWR.n521 VDPWR.n519 92.5005
R2596 VDPWR.n524 VDPWR.n521 92.5005
R2597 VDPWR.n520 VDPWR 92.5005
R2598 VDPWR.n522 VDPWR.n520 92.5005
R2599 VDPWR.n551 VDPWR.n528 92.5005
R2600 VDPWR.n528 VDPWR.n524 92.5005
R2601 VDPWR VDPWR.n527 92.5005
R2602 VDPWR.n527 VDPWR.n522 92.5005
R2603 VDPWR VDPWR.n539 92.5005
R2604 VDPWR.n539 VDPWR.n537 92.5005
R2605 VDPWR.n540 VDPWR.n538 92.5005
R2606 VDPWR.n538 VDPWR.n533 92.5005
R2607 VDPWR VDPWR.n30 92.5005
R2608 VDPWR.n30 VDPWR.n28 92.5005
R2609 VDPWR.n32 VDPWR.n29 92.5005
R2610 VDPWR.n29 VDPWR.n28 92.5005
R2611 VDPWR VDPWR.n15 92.5005
R2612 VDPWR.n15 VDPWR.n13 92.5005
R2613 VDPWR VDPWR.n70 92.5005
R2614 VDPWR.n70 VDPWR.n69 92.5005
R2615 VDPWR.n54 VDPWR 92.5005
R2616 VDPWR.n55 VDPWR.n54 92.5005
R2617 VDPWR.n57 VDPWR.n56 92.5005
R2618 VDPWR.n56 VDPWR.n55 92.5005
R2619 VDPWR.n68 VDPWR.n67 92.5005
R2620 VDPWR.n69 VDPWR.n68 92.5005
R2621 VDPWR.n16 VDPWR.n14 92.5005
R2622 VDPWR.n14 VDPWR.n13 92.5005
R2623 VDPWR VDPWR.n10 92.5005
R2624 VDPWR.n10 VDPWR.n8 92.5005
R2625 VDPWR.n12 VDPWR.n9 92.5005
R2626 VDPWR.n9 VDPWR.n8 92.5005
R2627 VDPWR.n83 VDPWR 92.5005
R2628 VDPWR.n5 VDPWR.n4 92.5005
R2629 VDPWR.n6 VDPWR.n5 92.5005
R2630 VDPWR VDPWR.n35 92.5005
R2631 VDPWR.n35 VDPWR.n33 92.5005
R2632 VDPWR.n40 VDPWR.n34 92.5005
R2633 VDPWR.n506 VDPWR.n474 91.6935
R2634 VDPWR.n506 VDPWR.n476 91.6935
R2635 VDPWR.n496 VDPWR.n485 91.6935
R2636 VDPWR.n496 VDPWR.n489 91.6935
R2637 VDPWR.n554 VDPWR.n522 91.6935
R2638 VDPWR.n554 VDPWR.n524 91.6935
R2639 VDPWR.n544 VDPWR.n533 91.6935
R2640 VDPWR.n544 VDPWR.n537 91.6935
R2641 VDPWR.n767 VDPWR.n752 89.559
R2642 VDPWR.n772 VDPWR.n752 89.559
R2643 VDPWR.n775 VDPWR.n748 89.559
R2644 VDPWR.n802 VDPWR.n748 89.559
R2645 VDPWR.n801 VDPWR.n780 89.559
R2646 VDPWR.n794 VDPWR.n780 89.559
R2647 VDPWR.n794 VDPWR.n793 89.559
R2648 VDPWR.n793 VDPWR.n787 89.559
R2649 VDPWR.n787 VDPWR.n739 89.559
R2650 VDPWR.n815 VDPWR.n739 89.559
R2651 VDPWR.n827 VDPWR.n816 89.559
R2652 VDPWR.n827 VDPWR.n722 89.559
R2653 VDPWR.n835 VDPWR.n722 89.559
R2654 VDPWR.n835 VDPWR.n672 89.559
R2655 VDPWR.n839 VDPWR.n672 89.559
R2656 VDPWR.n839 VDPWR.n716 89.559
R2657 VDPWR.n715 VDPWR.n675 89.559
R2658 VDPWR.n696 VDPWR.n675 89.559
R2659 VDPWR.n699 VDPWR.n685 89.559
R2660 VDPWR.n704 VDPWR.n685 89.559
R2661 VDPWR.n435 VDPWR.n330 85.0829
R2662 VDPWR.n436 VDPWR.n435 85.0829
R2663 VDPWR.n414 VDPWR.n375 85.0829
R2664 VDPWR.n390 VDPWR.n375 85.0829
R2665 VDPWR.n209 VDPWR.n188 85.0829
R2666 VDPWR.n209 VDPWR.n184 85.0829
R2667 VDPWR.n313 VDPWR.n312 85.0829
R2668 VDPWR.n312 VDPWR.n110 85.0829
R2669 VDPWR.n295 VDPWR.n98 85.0829
R2670 VDPWR.n296 VDPWR.n295 85.0829
R2671 VDPWR.n181 VDPWR.n175 85.0829
R2672 VDPWR.n175 VDPWR.n174 85.0829
R2673 VDPWR.n575 VDPWR.n574 85.0829
R2674 VDPWR.n574 VDPWR.n566 85.0829
R2675 VDPWR.n84 VDPWR.n83 79.4196
R2676 VDPWR.n41 VDPWR.n34 79.4196
R2677 VDPWR.n353 VDPWR.n341 66.7857
R2678 VDPWR.n397 VDPWR.n396 66.7857
R2679 VDPWR.n218 VDPWR.n217 66.7857
R2680 VDPWR.n141 VDPWR.n108 66.7857
R2681 VDPWR.n291 VDPWR.n131 66.7857
R2682 VDPWR.n238 VDPWR.n237 66.7857
R2683 VDPWR.n636 VDPWR.n635 66.7857
R2684 VDPWR.n431 VDPWR.n345 66.1931
R2685 VDPWR.n395 VDPWR.n394 66.1931
R2686 VDPWR.n216 VDPWR.n192 66.1931
R2687 VDPWR.n140 VDPWR.n117 66.1931
R2688 VDPWR.n130 VDPWR.n129 66.1931
R2689 VDPWR.n236 VDPWR.n235 66.1931
R2690 VDPWR.n590 VDPWR.n577 66.1931
R2691 VDPWR.n418 VDPWR.n417 62.6339
R2692 VDPWR.n445 VDPWR.n346 62.6339
R2693 VDPWR.n604 VDPWR.n587 62.6339
R2694 VDPWR.n256 VDPWR.n144 61.5478
R2695 VDPWR.n287 VDPWR.n137 61.5478
R2696 VDPWR.n201 VDPWR.n200 61.3667
R2697 VDPWR.n267 VDPWR.n122 61.3667
R2698 VDPWR.n403 VDPWR.n402 60.4616
R2699 VDPWR.n453 VDPWR.n452 60.4616
R2700 VDPWR.n639 VDPWR.n571 60.4616
R2701 VDPWR.n802 VDPWR.n801 60.084
R2702 VDPWR.n816 VDPWR.n815 60.084
R2703 VDPWR.n716 VDPWR.n715 60.084
R2704 VDPWR VDPWR.n720 59.4829
R2705 VDPWR VDPWR.n720 59.4829
R2706 VDPWR.n837 VDPWR 59.4829
R2707 VDPWR VDPWR.n837 59.4829
R2708 VDPWR.n824 VDPWR.n823 59.4829
R2709 VDPWR.n823 VDPWR.n667 59.4829
R2710 VDPWR.n842 VDPWR.n841 59.4829
R2711 VDPWR.n783 VDPWR 59.4829
R2712 VDPWR VDPWR.n783 59.4829
R2713 VDPWR VDPWR.n791 59.4829
R2714 VDPWR.n791 VDPWR 59.4829
R2715 VDPWR.n798 VDPWR.n797 59.4829
R2716 VDPWR.n797 VDPWR.n743 59.4829
R2717 VDPWR.n812 VDPWR.n811 59.4829
R2718 VDPWR.n832 VDPWR.n727 59.4829
R2719 VDPWR.n833 VDPWR.n832 59.4829
R2720 VDPWR.n732 VDPWR.n731 59.4829
R2721 VDPWR VDPWR.n736 59.4829
R2722 VDPWR.n736 VDPWR 59.4829
R2723 VDPWR VDPWR.n735 59.4829
R2724 VDPWR.n735 VDPWR 59.4829
R2725 VDPWR.n60 VDPWR.n57 59.4829
R2726 VDPWR.n67 VDPWR.n60 59.4829
R2727 VDPWR.n61 VDPWR.n16 59.4829
R2728 VDPWR VDPWR.n18 59.4829
R2729 VDPWR VDPWR.n18 59.4829
R2730 VDPWR.n71 VDPWR 59.4829
R2731 VDPWR VDPWR.n71 59.4829
R2732 VDPWR.n843 VDPWR.n842 59.1064
R2733 VDPWR.n811 VDPWR.n810 59.1064
R2734 VDPWR.n731 VDPWR.n665 59.1064
R2735 VDPWR.n66 VDPWR.n61 59.1064
R2736 VDPWR.n775 VDPWR.n772 58.9504
R2737 VDPWR.n699 VDPWR.n696 58.9504
R2738 VDPWR.n436 VDPWR.n432 52.3937
R2739 VDPWR.n390 VDPWR.n386 52.3937
R2740 VDPWR.n219 VDPWR.n188 52.3937
R2741 VDPWR.n314 VDPWR.n313 52.3937
R2742 VDPWR.n296 VDPWR.n292 52.3937
R2743 VDPWR.n174 VDPWR.n167 52.3937
R2744 VDPWR.n637 VDPWR.n575 52.3937
R2745 VDPWR.n438 VDPWR.n437 51.2005
R2746 VDPWR.n392 VDPWR.n391 51.2005
R2747 VDPWR.n205 VDPWR.n204 51.2005
R2748 VDPWR.n306 VDPWR.n109 51.2005
R2749 VDPWR.n298 VDPWR.n297 51.2005
R2750 VDPWR.n233 VDPWR.n170 51.2005
R2751 VDPWR.n602 VDPWR.n586 51.2005
R2752 VDPWR.n449 VDPWR.n448 37.0005
R2753 VDPWR.n448 VDPWR.n337 37.0005
R2754 VDPWR.n440 VDPWR.n344 37.0005
R2755 VDPWR.n426 VDPWR.n344 37.0005
R2756 VDPWR.n377 VDPWR.n376 37.0005
R2757 VDPWR.n377 VDPWR.n359 37.0005
R2758 VDPWR.n374 VDPWR.n372 37.0005
R2759 VDPWR.n372 VDPWR.n371 37.0005
R2760 VDPWR.n435 VDPWR.n434 37.0005
R2761 VDPWR.n434 VDPWR.n334 37.0005
R2762 VDPWR.n333 VDPWR.n331 37.0005
R2763 VDPWR.n339 VDPWR.n333 37.0005
R2764 VDPWR.n442 VDPWR.n348 37.0005
R2765 VDPWR.n427 VDPWR.n348 37.0005
R2766 VDPWR.n400 VDPWR.n399 37.0005
R2767 VDPWR.n401 VDPWR.n400 37.0005
R2768 VDPWR.n389 VDPWR.n388 37.0005
R2769 VDPWR.n388 VDPWR.n367 37.0005
R2770 VDPWR.n381 VDPWR.n375 37.0005
R2771 VDPWR.n381 VDPWR.n380 37.0005
R2772 VDPWR.n280 VDPWR.n132 37.0005
R2773 VDPWR.n281 VDPWR.n280 37.0005
R2774 VDPWR.n301 VDPWR.n300 37.0005
R2775 VDPWR.n302 VDPWR.n301 37.0005
R2776 VDPWR.n229 VDPWR.n228 37.0005
R2777 VDPWR.n229 VDPWR.n144 37.0005
R2778 VDPWR.n177 VDPWR.n171 37.0005
R2779 VDPWR.n201 VDPWR.n171 37.0005
R2780 VDPWR.n295 VDPWR.n294 37.0005
R2781 VDPWR.n294 VDPWR.n102 37.0005
R2782 VDPWR.n101 VDPWR.n99 37.0005
R2783 VDPWR.n137 VDPWR.n101 37.0005
R2784 VDPWR.n127 VDPWR.n126 37.0005
R2785 VDPWR.n126 VDPWR.n122 37.0005
R2786 VDPWR.n210 VDPWR.n209 37.0005
R2787 VDPWR.n213 VDPWR.n210 37.0005
R2788 VDPWR.n221 VDPWR.n185 37.0005
R2789 VDPWR.n221 VDPWR.n144 37.0005
R2790 VDPWR.n202 VDPWR.n199 37.0005
R2791 VDPWR.n202 VDPWR.n201 37.0005
R2792 VDPWR.n312 VDPWR.n311 37.0005
R2793 VDPWR.n311 VDPWR.n102 37.0005
R2794 VDPWR.n278 VDPWR.n107 37.0005
R2795 VDPWR.n137 VDPWR.n107 37.0005
R2796 VDPWR.n118 VDPWR.n111 37.0005
R2797 VDPWR.n122 VDPWR.n111 37.0005
R2798 VDPWR.n190 VDPWR.n164 37.0005
R2799 VDPWR.n242 VDPWR.n164 37.0005
R2800 VDPWR.n196 VDPWR.n193 37.0005
R2801 VDPWR.n193 VDPWR.n153 37.0005
R2802 VDPWR.n283 VDPWR.n282 37.0005
R2803 VDPWR.n282 VDPWR.n281 37.0005
R2804 VDPWR.n304 VDPWR.n303 37.0005
R2805 VDPWR.n303 VDPWR.n302 37.0005
R2806 VDPWR.n241 VDPWR.n240 37.0005
R2807 VDPWR.n242 VDPWR.n241 37.0005
R2808 VDPWR.n169 VDPWR.n168 37.0005
R2809 VDPWR.n168 VDPWR.n153 37.0005
R2810 VDPWR.n175 VDPWR.n172 37.0005
R2811 VDPWR.n213 VDPWR.n172 37.0005
R2812 VDPWR.n574 VDPWR.n573 37.0005
R2813 VDPWR.n573 VDPWR.n570 37.0005
R2814 VDPWR.n569 VDPWR.n567 37.0005
R2815 VDPWR.n611 VDPWR.n569 37.0005
R2816 VDPWR.n598 VDPWR.n589 37.0005
R2817 VDPWR.n594 VDPWR.n589 37.0005
R2818 VDPWR.n609 VDPWR.n608 37.0005
R2819 VDPWR.n610 VDPWR.n609 37.0005
R2820 VDPWR.n600 VDPWR.n585 37.0005
R2821 VDPWR.n593 VDPWR.n585 37.0005
R2822 VDPWR VDPWR.n618 37.0005
R2823 VDPWR.n627 VDPWR.n626 37.0005
R2824 VDPWR.n628 VDPWR.n627 37.0005
R2825 VDPWR.n249 VDPWR.n156 31.3172
R2826 VDPWR.n308 VDPWR.n113 31.3172
R2827 VDPWR.n243 VDPWR.n162 30.2311
R2828 VDPWR.n316 VDPWR.n105 30.2311
R2829 VDPWR.n441 VDPWR.n349 26.6787
R2830 VDPWR.n387 VDPWR.n364 26.6787
R2831 VDPWR.n197 VDPWR.n159 26.6787
R2832 VDPWR.n143 VDPWR.n119 26.6787
R2833 VDPWR.n265 VDPWR.n128 26.6787
R2834 VDPWR.n176 VDPWR.n150 26.6787
R2835 VDPWR.n599 VDPWR.n596 26.6787
R2836 VDPWR.n351 VDPWR.n342 26.63
R2837 VDPWR.n423 VDPWR.n362 26.63
R2838 VDPWR.n189 VDPWR.n161 26.63
R2839 VDPWR.n285 VDPWR.n284 26.63
R2840 VDPWR.n136 VDPWR.n135 26.63
R2841 VDPWR.n254 VDPWR.n148 26.63
R2842 VDPWR.n607 VDPWR.n583 26.63
R2843 VDPWR.n485 VDPWR.n476 26.5564
R2844 VDPWR.n533 VDPWR.n524 26.5564
R2845 VDPWR.n779 VDPWR.n778 23.1255
R2846 VDPWR.n802 VDPWR.n779 23.1255
R2847 VDPWR.n777 VDPWR.n776 23.1255
R2848 VDPWR.n776 VDPWR.n775 23.1255
R2849 VDPWR.n831 VDPWR.n830 23.1255
R2850 VDPWR.n830 VDPWR.n722 23.1255
R2851 VDPWR.n730 VDPWR.n729 23.1255
R2852 VDPWR.n729 VDPWR.n672 23.1255
R2853 VDPWR.n734 VDPWR.n733 23.1255
R2854 VDPWR.n733 VDPWR.n716 23.1255
R2855 VDPWR.n738 VDPWR.n737 23.1255
R2856 VDPWR.n816 VDPWR.n737 23.1255
R2857 VDPWR.n694 VDPWR.n693 23.1255
R2858 VDPWR.n696 VDPWR.n694 23.1255
R2859 VDPWR.n692 VDPWR.n674 23.1255
R2860 VDPWR.n715 VDPWR.n674 23.1255
R2861 VDPWR.n703 VDPWR.n702 23.1255
R2862 VDPWR.n704 VDPWR.n703 23.1255
R2863 VDPWR.n701 VDPWR.n700 23.1255
R2864 VDPWR.n700 VDPWR.n699 23.1255
R2865 VDPWR.n760 VDPWR.n753 23.1255
R2866 VDPWR.n772 VDPWR.n753 23.1255
R2867 VDPWR.n766 VDPWR.n765 23.1255
R2868 VDPWR.n767 VDPWR.n766 23.1255
R2869 VDPWR.n804 VDPWR.n803 23.1255
R2870 VDPWR.n803 VDPWR.n802 23.1255
R2871 VDPWR.n774 VDPWR.n773 23.1255
R2872 VDPWR.n775 VDPWR.n774 23.1255
R2873 VDPWR.n796 VDPWR.n795 23.1255
R2874 VDPWR.n795 VDPWR.n794 23.1255
R2875 VDPWR.n789 VDPWR.n742 23.1255
R2876 VDPWR.n789 VDPWR.n787 23.1255
R2877 VDPWR.n814 VDPWR.n813 23.1255
R2878 VDPWR.n815 VDPWR.n814 23.1255
R2879 VDPWR.n800 VDPWR.n799 23.1255
R2880 VDPWR.n801 VDPWR.n800 23.1255
R2881 VDPWR.n822 VDPWR.n821 23.1255
R2882 VDPWR.n821 VDPWR.n722 23.1255
R2883 VDPWR.n718 VDPWR.n668 23.1255
R2884 VDPWR.n718 VDPWR.n672 23.1255
R2885 VDPWR.n671 VDPWR.n669 23.1255
R2886 VDPWR.n716 VDPWR.n671 23.1255
R2887 VDPWR.n825 VDPWR.n819 23.1255
R2888 VDPWR.n819 VDPWR.n816 23.1255
R2889 VDPWR.n695 VDPWR.n678 23.1255
R2890 VDPWR.n696 VDPWR.n695 23.1255
R2891 VDPWR.n714 VDPWR.n713 23.1255
R2892 VDPWR.n715 VDPWR.n714 23.1255
R2893 VDPWR.n706 VDPWR.n705 23.1255
R2894 VDPWR.n705 VDPWR.n704 23.1255
R2895 VDPWR.n698 VDPWR.n697 23.1255
R2896 VDPWR.n699 VDPWR.n698 23.1255
R2897 VDPWR.n771 VDPWR.n770 23.1255
R2898 VDPWR.n772 VDPWR.n771 23.1255
R2899 VDPWR.n769 VDPWR.n768 23.1255
R2900 VDPWR.n768 VDPWR.n767 23.1255
R2901 VDPWR.n498 VDPWR.n497 23.1255
R2902 VDPWR.n497 VDPWR.n496 23.1255
R2903 VDPWR.n488 VDPWR.n487 23.1255
R2904 VDPWR.n496 VDPWR.n488 23.1255
R2905 VDPWR.n508 VDPWR.n507 23.1255
R2906 VDPWR.n507 VDPWR.n506 23.1255
R2907 VDPWR.n478 VDPWR.n477 23.1255
R2908 VDPWR.n506 VDPWR.n478 23.1255
R2909 VDPWR.n481 VDPWR.n475 23.1255
R2910 VDPWR.n506 VDPWR.n475 23.1255
R2911 VDPWR.n505 VDPWR.n504 23.1255
R2912 VDPWR.n506 VDPWR.n505 23.1255
R2913 VDPWR.n495 VDPWR.n494 23.1255
R2914 VDPWR.n496 VDPWR.n495 23.1255
R2915 VDPWR.n493 VDPWR.n486 23.1255
R2916 VDPWR.n496 VDPWR.n486 23.1255
R2917 VDPWR.n546 VDPWR.n545 23.1255
R2918 VDPWR.n545 VDPWR.n544 23.1255
R2919 VDPWR.n536 VDPWR.n535 23.1255
R2920 VDPWR.n544 VDPWR.n536 23.1255
R2921 VDPWR.n556 VDPWR.n555 23.1255
R2922 VDPWR.n555 VDPWR.n554 23.1255
R2923 VDPWR.n526 VDPWR.n525 23.1255
R2924 VDPWR.n554 VDPWR.n526 23.1255
R2925 VDPWR.n529 VDPWR.n523 23.1255
R2926 VDPWR.n554 VDPWR.n523 23.1255
R2927 VDPWR.n553 VDPWR.n552 23.1255
R2928 VDPWR.n554 VDPWR.n553 23.1255
R2929 VDPWR.n543 VDPWR.n542 23.1255
R2930 VDPWR.n544 VDPWR.n543 23.1255
R2931 VDPWR.n541 VDPWR.n534 23.1255
R2932 VDPWR.n544 VDPWR.n534 23.1255
R2933 VDPWR.n51 VDPWR.n50 23.1255
R2934 VDPWR.n52 VDPWR.n51 23.1255
R2935 VDPWR.n49 VDPWR.n48 23.1255
R2936 VDPWR.n48 VDPWR.n47 23.1255
R2937 VDPWR.n59 VDPWR.n58 23.1255
R2938 VDPWR.n58 VDPWR.n21 23.1255
R2939 VDPWR.n24 VDPWR.n17 23.1255
R2940 VDPWR.n24 VDPWR.n22 23.1255
R2941 VDPWR.n73 VDPWR.n72 23.1255
R2942 VDPWR.n74 VDPWR.n73 23.1255
R2943 VDPWR.n27 VDPWR.n26 23.1255
R2944 VDPWR.n53 VDPWR.n27 23.1255
R2945 VDPWR.n79 VDPWR.n78 23.1255
R2946 VDPWR.n80 VDPWR.n79 23.1255
R2947 VDPWR.n77 VDPWR.n76 23.1255
R2948 VDPWR.n76 VDPWR.n75 23.1255
R2949 VDPWR.n86 VDPWR.n85 23.1255
R2950 VDPWR.n82 VDPWR.n7 23.1255
R2951 VDPWR.n82 VDPWR.n81 23.1255
R2952 VDPWR.n45 VDPWR.n44 23.1255
R2953 VDPWR.n46 VDPWR.n45 23.1255
R2954 VDPWR.n43 VDPWR.n42 23.1255
R2955 VDPWR.n439 VDPWR.n438 19.0689
R2956 VDPWR.n393 VDPWR.n392 19.0689
R2957 VDPWR.n204 VDPWR.n194 19.0689
R2958 VDPWR.n306 VDPWR.n305 19.0689
R2959 VDPWR.n299 VDPWR.n298 19.0689
R2960 VDPWR.n234 VDPWR.n233 19.0689
R2961 VDPWR.n602 VDPWR.n601 19.0689
R2962 VDPWR.n418 VDPWR.n367 17.7406
R2963 VDPWR.n426 VDPWR.n346 17.7406
R2964 VDPWR.n593 VDPWR.n587 17.7406
R2965 VDPWR.n449 VDPWR.n342 17.4344
R2966 VDPWR.n399 VDPWR.n362 17.4344
R2967 VDPWR.n190 VDPWR.n189 17.4344
R2968 VDPWR.n284 VDPWR.n283 17.4344
R2969 VDPWR.n135 VDPWR.n132 17.4344
R2970 VDPWR.n240 VDPWR.n148 17.4344
R2971 VDPWR.n608 VDPWR.n607 17.4344
R2972 VDPWR.n397 VDPWR.n386 16.8923
R2973 VDPWR.n432 VDPWR.n341 16.8923
R2974 VDPWR.n238 VDPWR.n167 16.8923
R2975 VDPWR.n219 VDPWR.n218 16.8923
R2976 VDPWR.n314 VDPWR.n108 16.8923
R2977 VDPWR.n292 VDPWR.n291 16.8923
R2978 VDPWR.n637 VDPWR.n636 16.8923
R2979 VDPWR.n441 VDPWR.n440 16.6793
R2980 VDPWR.n389 VDPWR.n387 16.6793
R2981 VDPWR.n197 VDPWR.n196 16.6793
R2982 VDPWR.n304 VDPWR.n119 16.6793
R2983 VDPWR.n300 VDPWR.n128 16.6793
R2984 VDPWR.n176 VDPWR.n169 16.6793
R2985 VDPWR.n600 VDPWR.n599 16.6793
R2986 VDPWR.n355 VDPWR.n354 14.2313
R2987 VDPWR.n354 VDPWR.n334 14.2313
R2988 VDPWR.n351 VDPWR.n340 14.2313
R2989 VDPWR.n429 VDPWR.n349 14.2313
R2990 VDPWR.n429 VDPWR.n428 14.2313
R2991 VDPWR.n424 VDPWR.n423 14.2313
R2992 VDPWR.n425 VDPWR.n424 14.2313
R2993 VDPWR.n379 VDPWR.n363 14.2313
R2994 VDPWR.n380 VDPWR.n379 14.2313
R2995 VDPWR.n365 VDPWR.n364 14.2313
R2996 VDPWR.n262 VDPWR.n261 14.2313
R2997 VDPWR.n261 VDPWR.n102 14.2313
R2998 VDPWR.n288 VDPWR.n136 14.2313
R2999 VDPWR.n288 VDPWR.n287 14.2313
R3000 VDPWR.n266 VDPWR.n265 14.2313
R3001 VDPWR.n267 VDPWR.n266 14.2313
R3002 VDPWR.n212 VDPWR.n160 14.2313
R3003 VDPWR.n213 VDPWR.n212 14.2313
R3004 VDPWR.n161 VDPWR.n145 14.2313
R3005 VDPWR.n256 VDPWR.n145 14.2313
R3006 VDPWR.n159 VDPWR.n157 14.2313
R3007 VDPWR.n200 VDPWR.n157 14.2313
R3008 VDPWR.n271 VDPWR.n142 14.2313
R3009 VDPWR.n271 VDPWR.n102 14.2313
R3010 VDPWR.n286 VDPWR.n285 14.2313
R3011 VDPWR.n287 VDPWR.n286 14.2313
R3012 VDPWR.n268 VDPWR.n143 14.2313
R3013 VDPWR.n268 VDPWR.n267 14.2313
R3014 VDPWR.n255 VDPWR.n254 14.2313
R3015 VDPWR.n256 VDPWR.n255 14.2313
R3016 VDPWR.n208 VDPWR.n149 14.2313
R3017 VDPWR.n213 VDPWR.n208 14.2313
R3018 VDPWR.n151 VDPWR.n150 14.2313
R3019 VDPWR.n200 VDPWR.n151 14.2313
R3020 VDPWR.n634 VDPWR.n633 14.2313
R3021 VDPWR.n633 VDPWR.n570 14.2313
R3022 VDPWR.n630 VDPWR.n583 14.2313
R3023 VDPWR.n630 VDPWR.n629 14.2313
R3024 VDPWR.n596 VDPWR.n595 14.2313
R3025 VDPWR.n84 VDPWR.n6 8.97701
R3026 VDPWR.n41 VDPWR.n33 8.97701
R3027 VDPWR.n249 VDPWR.n153 8.87055
R3028 VDPWR.n302 VDPWR.n113 8.87055
R3029 VDPWR.n380 VDPWR.n370 7.96544
R3030 VDPWR.n446 VDPWR.n334 7.96544
R3031 VDPWR.n605 VDPWR.n570 7.96544
R3032 VDPWR.n432 VDPWR.n335 7.11588
R3033 VDPWR.n453 VDPWR.n335 7.11588
R3034 VDPWR.n438 VDPWR.n347 7.11588
R3035 VDPWR.n445 VDPWR.n347 7.11588
R3036 VDPWR.n444 VDPWR.n443 7.11588
R3037 VDPWR.n445 VDPWR.n444 7.11588
R3038 VDPWR.n455 VDPWR.n454 7.11588
R3039 VDPWR.n454 VDPWR.n453 7.11588
R3040 VDPWR.n386 VDPWR.n383 7.11588
R3041 VDPWR.n403 VDPWR.n383 7.11588
R3042 VDPWR.n392 VDPWR.n369 7.11588
R3043 VDPWR.n417 VDPWR.n369 7.11588
R3044 VDPWR.n416 VDPWR.n415 7.11588
R3045 VDPWR.n417 VDPWR.n416 7.11588
R3046 VDPWR.n405 VDPWR.n404 7.11588
R3047 VDPWR.n404 VDPWR.n403 7.11588
R3048 VDPWR.n292 VDPWR.n104 7.11588
R3049 VDPWR.n316 VDPWR.n104 7.11588
R3050 VDPWR.n298 VDPWR.n114 7.11588
R3051 VDPWR.n308 VDPWR.n114 7.11588
R3052 VDPWR.n125 VDPWR.n116 7.11588
R3053 VDPWR.n308 VDPWR.n116 7.11588
R3054 VDPWR.n318 VDPWR.n317 7.11588
R3055 VDPWR.n317 VDPWR.n316 7.11588
R3056 VDPWR.n223 VDPWR.n222 7.11588
R3057 VDPWR.n222 VDPWR.n162 7.11588
R3058 VDPWR.n198 VDPWR.n195 7.11588
R3059 VDPWR.n195 VDPWR.n156 7.11588
R3060 VDPWR.n204 VDPWR.n203 7.11588
R3061 VDPWR.n203 VDPWR.n156 7.11588
R3062 VDPWR.n220 VDPWR.n219 7.11588
R3063 VDPWR.n220 VDPWR.n162 7.11588
R3064 VDPWR.n277 VDPWR.n103 7.11588
R3065 VDPWR.n316 VDPWR.n103 7.11588
R3066 VDPWR.n309 VDPWR.n112 7.11588
R3067 VDPWR.n309 VDPWR.n308 7.11588
R3068 VDPWR.n307 VDPWR.n306 7.11588
R3069 VDPWR.n308 VDPWR.n307 7.11588
R3070 VDPWR.n315 VDPWR.n314 7.11588
R3071 VDPWR.n316 VDPWR.n315 7.11588
R3072 VDPWR.n230 VDPWR.n167 7.11588
R3073 VDPWR.n230 VDPWR.n162 7.11588
R3074 VDPWR.n233 VDPWR.n232 7.11588
R3075 VDPWR.n232 VDPWR.n156 7.11588
R3076 VDPWR.n180 VDPWR.n179 7.11588
R3077 VDPWR.n179 VDPWR.n156 7.11588
R3078 VDPWR.n227 VDPWR.n173 7.11588
R3079 VDPWR.n173 VDPWR.n162 7.11588
R3080 VDPWR.n641 VDPWR.n640 7.11588
R3081 VDPWR.n640 VDPWR.n639 7.11588
R3082 VDPWR.n597 VDPWR.n588 7.11588
R3083 VDPWR.n604 VDPWR.n588 7.11588
R3084 VDPWR.n603 VDPWR.n602 7.11588
R3085 VDPWR.n604 VDPWR.n603 7.11588
R3086 VDPWR.n638 VDPWR.n637 7.11588
R3087 VDPWR.n639 VDPWR.n638 7.11588
R3088 VDPWR.n323 VDPWR 6.74008
R3089 VDPWR.n460 VDPWR 6.737
R3090 VDPWR.n323 VDPWR 6.73352
R3091 VDPWR.n409 VDPWR.n408 6.63939
R3092 VDPWR.n647 VDPWR.n646 6.63939
R3093 VDPWR.n352 VDPWR.n336 5.78175
R3094 VDPWR.n452 VDPWR.n336 5.78175
R3095 VDPWR.n358 VDPWR.n357 5.78175
R3096 VDPWR.n358 VDPWR.n346 5.78175
R3097 VDPWR.n431 VDPWR.n430 5.78175
R3098 VDPWR.n430 VDPWR.n346 5.78175
R3099 VDPWR.n451 VDPWR.n450 5.78175
R3100 VDPWR.n452 VDPWR.n451 5.78175
R3101 VDPWR.n447 VDPWR.n345 5.78175
R3102 VDPWR.n447 VDPWR.n446 5.78175
R3103 VDPWR.n437 VDPWR.n343 5.78175
R3104 VDPWR.n446 VDPWR.n343 5.78175
R3105 VDPWR.n398 VDPWR.n360 5.78175
R3106 VDPWR.n402 VDPWR.n360 5.78175
R3107 VDPWR.n394 VDPWR.n368 5.78175
R3108 VDPWR.n418 VDPWR.n368 5.78175
R3109 VDPWR.n395 VDPWR.n385 5.78175
R3110 VDPWR.n385 VDPWR.n370 5.78175
R3111 VDPWR.n422 VDPWR.n361 5.78175
R3112 VDPWR.n402 VDPWR.n361 5.78175
R3113 VDPWR.n420 VDPWR.n419 5.78175
R3114 VDPWR.n419 VDPWR.n418 5.78175
R3115 VDPWR.n391 VDPWR.n384 5.78175
R3116 VDPWR.n384 VDPWR.n370 5.78175
R3117 VDPWR.n259 VDPWR.n134 5.78175
R3118 VDPWR.n134 VDPWR.n105 5.78175
R3119 VDPWR.n264 VDPWR.n258 5.78175
R3120 VDPWR.n258 VDPWR.n113 5.78175
R3121 VDPWR.n257 VDPWR.n129 5.78175
R3122 VDPWR.n257 VDPWR.n113 5.78175
R3123 VDPWR.n290 VDPWR.n289 5.78175
R3124 VDPWR.n289 VDPWR.n105 5.78175
R3125 VDPWR.n130 VDPWR.n124 5.78175
R3126 VDPWR.n124 VDPWR.n115 5.78175
R3127 VDPWR.n297 VDPWR.n123 5.78175
R3128 VDPWR.n123 VDPWR.n115 5.78175
R3129 VDPWR.n206 VDPWR.n205 5.78175
R3130 VDPWR.n214 VDPWR.n206 5.78175
R3131 VDPWR.n216 VDPWR.n215 5.78175
R3132 VDPWR.n215 VDPWR.n214 5.78175
R3133 VDPWR.n121 VDPWR.n109 5.78175
R3134 VDPWR.n121 VDPWR.n115 5.78175
R3135 VDPWR.n140 VDPWR.n120 5.78175
R3136 VDPWR.n120 VDPWR.n115 5.78175
R3137 VDPWR.n191 VDPWR.n163 5.78175
R3138 VDPWR.n243 VDPWR.n163 5.78175
R3139 VDPWR.n192 VDPWR.n155 5.78175
R3140 VDPWR.n249 VDPWR.n155 5.78175
R3141 VDPWR.n248 VDPWR.n247 5.78175
R3142 VDPWR.n249 VDPWR.n248 5.78175
R3143 VDPWR.n245 VDPWR.n244 5.78175
R3144 VDPWR.n244 VDPWR.n243 5.78175
R3145 VDPWR.n279 VDPWR.n139 5.78175
R3146 VDPWR.n139 VDPWR.n105 5.78175
R3147 VDPWR.n269 VDPWR.n117 5.78175
R3148 VDPWR.n269 VDPWR.n113 5.78175
R3149 VDPWR.n274 VDPWR.n273 5.78175
R3150 VDPWR.n273 VDPWR.n113 5.78175
R3151 VDPWR.n276 VDPWR.n138 5.78175
R3152 VDPWR.n138 VDPWR.n105 5.78175
R3153 VDPWR.n239 VDPWR.n146 5.78175
R3154 VDPWR.n243 VDPWR.n146 5.78175
R3155 VDPWR.n235 VDPWR.n154 5.78175
R3156 VDPWR.n249 VDPWR.n154 5.78175
R3157 VDPWR.n236 VDPWR.n166 5.78175
R3158 VDPWR.n214 VDPWR.n166 5.78175
R3159 VDPWR.n253 VDPWR.n147 5.78175
R3160 VDPWR.n243 VDPWR.n147 5.78175
R3161 VDPWR.n251 VDPWR.n250 5.78175
R3162 VDPWR.n250 VDPWR.n249 5.78175
R3163 VDPWR.n170 VDPWR.n165 5.78175
R3164 VDPWR.n214 VDPWR.n165 5.78175
R3165 VDPWR.n606 VDPWR.n586 5.78175
R3166 VDPWR.n606 VDPWR.n605 5.78175
R3167 VDPWR.n584 VDPWR.n577 5.78175
R3168 VDPWR.n605 VDPWR.n584 5.78175
R3169 VDPWR.n631 VDPWR.n576 5.78175
R3170 VDPWR.n631 VDPWR.n571 5.78175
R3171 VDPWR.n590 VDPWR.n580 5.78175
R3172 VDPWR.n587 VDPWR.n580 5.78175
R3173 VDPWR.n592 VDPWR.n591 5.78175
R3174 VDPWR.n592 VDPWR.n587 5.78175
R3175 VDPWR.n582 VDPWR.n581 5.78175
R3176 VDPWR.n581 VDPWR.n571 5.78175
R3177 VDPWR.n615 VDPWR.n613 5.78175
R3178 VDPWR.n620 VDPWR.n614 5.78175
R3179 VDPWR.n614 VDPWR.n612 5.78175
R3180 VDPWR.n625 VDPWR.n620 4.71629
R3181 VDPWR.n376 VDPWR.n362 4.7119
R3182 VDPWR.n342 VDPWR.n331 4.7119
R3183 VDPWR.n189 VDPWR.n185 4.7119
R3184 VDPWR.n228 VDPWR.n148 4.7119
R3185 VDPWR.n284 VDPWR.n278 4.7119
R3186 VDPWR.n135 VDPWR.n99 4.7119
R3187 VDPWR.n607 VDPWR.n567 4.7119
R3188 VDPWR.n387 VDPWR.n374 4.70083
R3189 VDPWR.n442 VDPWR.n441 4.70083
R3190 VDPWR.n199 VDPWR.n197 4.70083
R3191 VDPWR.n177 VDPWR.n176 4.70083
R3192 VDPWR.n119 VDPWR.n118 4.70083
R3193 VDPWR.n128 VDPWR.n127 4.70083
R3194 VDPWR.n599 VDPWR.n598 4.70083
R3195 VDPWR.n617 VDPWR.n613 4.37746
R3196 VDPWR.n402 VDPWR.n401 3.98297
R3197 VDPWR.n452 VDPWR.n337 3.98297
R3198 VDPWR.n214 VDPWR.n213 3.98297
R3199 VDPWR.n115 VDPWR.n102 3.98297
R3200 VDPWR.n610 VDPWR.n571 3.98297
R3201 VDPWR.n652 VDPWR 3.64817
R3202 VDPWR.n322 VDPWR 3.52106
R3203 VDPWR.n92 VDPWR 3.52106
R3204 VDPWR.n659 VDPWR.n658 3.32168
R3205 VDPWR VDPWR.n0 3.05185
R3206 VDPWR.n563 VDPWR 2.62366
R3207 VDPWR.n761 VDPWR 2.3405
R3208 VDPWR.n761 VDPWR 2.3405
R3209 VDPWR.n807 VDPWR 2.3405
R3210 VDPWR.n807 VDPWR 2.3405
R3211 VDPWR.n709 VDPWR 2.3405
R3212 VDPWR.n709 VDPWR 2.3405
R3213 VDPWR.n681 VDPWR 2.3405
R3214 VDPWR.n681 VDPWR 2.3405
R3215 VDPWR.n470 VDPWR 2.3405
R3216 VDPWR.n470 VDPWR 2.3405
R3217 VDPWR.n500 VDPWR 2.3405
R3218 VDPWR.n500 VDPWR 2.3405
R3219 VDPWR.n518 VDPWR 2.3405
R3220 VDPWR.n518 VDPWR 2.3405
R3221 VDPWR.n548 VDPWR 2.3405
R3222 VDPWR.n548 VDPWR 2.3405
R3223 VDPWR.n89 VDPWR 2.3405
R3224 VDPWR.n62 VDPWR 2.3405
R3225 VDPWR.n36 VDPWR 2.3405
R3226 VDPWR.n38 VDPWR 2.3405
R3227 VDPWR.n808 VDPWR 2.29412
R3228 VDPWR.n666 VDPWR 2.29412
R3229 VDPWR.n666 VDPWR 2.29412
R3230 VDPWR.n64 VDPWR 2.29412
R3231 VDPWR.n243 VDPWR.n242 1.99173
R3232 VDPWR.n281 VDPWR.n105 1.99173
R3233 VDPWR.n97 VDPWR 1.93224
R3234 VDPWR.n183 VDPWR 1.93224
R3235 VDPWR.n39 VDPWR.n38 1.92169
R3236 VDPWR.n459 VDPWR 1.89811
R3237 VDPWR.n407 VDPWR 1.89811
R3238 VDPWR.n762 VDPWR.n756 1.8605
R3239 VDPWR.n806 VDPWR.n744 1.8605
R3240 VDPWR.n710 VDPWR.n679 1.8605
R3241 VDPWR.n708 VDPWR.n680 1.8605
R3242 VDPWR.n763 VDPWR.n762 1.8605
R3243 VDPWR.n806 VDPWR.n805 1.8605
R3244 VDPWR.n711 VDPWR.n710 1.8605
R3245 VDPWR.n708 VDPWR.n707 1.8605
R3246 VDPWR.n510 VDPWR.n469 1.8605
R3247 VDPWR.n501 VDPWR.n499 1.8605
R3248 VDPWR.n510 VDPWR.n509 1.8605
R3249 VDPWR.n502 VDPWR.n501 1.8605
R3250 VDPWR.n558 VDPWR.n517 1.8605
R3251 VDPWR.n549 VDPWR.n547 1.8605
R3252 VDPWR.n558 VDPWR.n557 1.8605
R3253 VDPWR.n550 VDPWR.n549 1.8605
R3254 VDPWR.n37 VDPWR.n31 1.8605
R3255 VDPWR.n63 VDPWR.n11 1.8605
R3256 VDPWR.n88 VDPWR.n87 1.8605
R3257 VDPWR.n439 VDPWR.n431 1.77828
R3258 VDPWR.n394 VDPWR.n393 1.77828
R3259 VDPWR.n194 VDPWR.n192 1.77828
R3260 VDPWR.n305 VDPWR.n117 1.77828
R3261 VDPWR.n299 VDPWR.n129 1.77828
R3262 VDPWR.n235 VDPWR.n234 1.77828
R3263 VDPWR.n601 VDPWR.n590 1.77828
R3264 VDPWR.n847 VDPWR.n846 1.76063
R3265 VDPWR.n560 VDPWR.n559 1.76063
R3266 VDPWR.n464 VDPWR.n324 1.753
R3267 VDPWR.n657 VDPWR.n656 1.753
R3268 VDPWR.n512 VDPWR.n511 1.75125
R3269 VDPWR.n326 VDPWR.n325 1.603
R3270 VDPWR.n462 VDPWR.n461 1.603
R3271 VDPWR.n644 VDPWR 1.43984
R3272 VDPWR.n617 VDPWR.n612 1.40064
R3273 VDPWR.n353 VDPWR.n345 1.3042
R3274 VDPWR.n396 VDPWR.n395 1.3042
R3275 VDPWR.n217 VDPWR.n216 1.3042
R3276 VDPWR.n141 VDPWR.n140 1.3042
R3277 VDPWR.n131 VDPWR.n130 1.3042
R3278 VDPWR.n237 VDPWR.n236 1.3042
R3279 VDPWR.n635 VDPWR.n577 1.3042
R3280 VDPWR.n437 VDPWR.n436 1.19372
R3281 VDPWR.n391 VDPWR.n390 1.19372
R3282 VDPWR.n205 VDPWR.n188 1.19372
R3283 VDPWR.n313 VDPWR.n109 1.19372
R3284 VDPWR.n297 VDPWR.n296 1.19372
R3285 VDPWR.n174 VDPWR.n170 1.19372
R3286 VDPWR.n586 VDPWR.n575 1.19372
R3287 VDPWR.n653 VDPWR.n3 1.18677
R3288 VDPWR.n846 VDPWR.n664 1.12394
R3289 VDPWR.n564 VDPWR.n465 1.10237
R3290 VDPWR.n511 VDPWR.n2 1.06531
R3291 VDPWR.n565 VDPWR 1.06379
R3292 VDPWR.n511 VDPWR.n510 1.06168
R3293 VDPWR.n559 VDPWR.n558 1.06168
R3294 VDPWR.n559 VDPWR.n516 1.05594
R3295 VDPWR.n329 VDPWR 1.04172
R3296 VDPWR.n411 VDPWR 1.04172
R3297 VDPWR.n321 VDPWR 0.890303
R3298 VDPWR.n182 VDPWR 0.890303
R3299 VDPWR.n621 VDPWR 0.85529
R3300 VDPWR.n458 VDPWR 0.854351
R3301 VDPWR.n406 VDPWR 0.854351
R3302 VDPWR.n562 VDPWR.n468 0.770146
R3303 VDPWR.n647 VDPWR 0.768852
R3304 VDPWR.n649 VDPWR.n648 0.73918
R3305 VDPWR.n844 VDPWR.n665 0.715885
R3306 VDPWR.n810 VDPWR.n809 0.715885
R3307 VDPWR.n844 VDPWR.n843 0.715885
R3308 VDPWR.n66 VDPWR.n65 0.715885
R3309 VDPWR.n408 VDPWR 0.69425
R3310 VDPWR.n460 VDPWR 0.69425
R3311 VDPWR.n562 VDPWR.n561 0.623777
R3312 VDPWR.n645 VDPWR.n644 0.619997
R3313 VDPWR.n565 VDPWR.n563 0.619997
R3314 VDPWR.n661 VDPWR.n90 0.615521
R3315 VDPWR.n90 VDPWR 0.559955
R3316 VDPWR.n97 VDPWR.n96 0.518921
R3317 VDPWR.n322 VDPWR.n321 0.518921
R3318 VDPWR.n183 VDPWR.n93 0.518921
R3319 VDPWR.n182 VDPWR.n92 0.518921
R3320 VDPWR.n652 VDPWR.n651 0.507812
R3321 VDPWR.n654 VDPWR.n653 0.507416
R3322 VDPWR.n95 VDPWR 0.505434
R3323 VDPWR.n658 VDPWR 0.505434
R3324 VDPWR.n329 VDPWR.n328 0.497975
R3325 VDPWR.n459 VDPWR.n458 0.497975
R3326 VDPWR.n407 VDPWR.n406 0.497975
R3327 VDPWR.n411 VDPWR.n410 0.497975
R3328 VDPWR.n659 VDPWR 0.467672
R3329 VDPWR.n323 VDPWR 0.467461
R3330 VDPWR VDPWR.n0 0.464224
R3331 VDPWR.n660 VDPWR.n659 0.426664
R3332 VDPWR.n809 VDPWR 0.413
R3333 VDPWR.n845 VDPWR.n844 0.410656
R3334 VDPWR.n707 VDPWR.n682 0.376971
R3335 VDPWR.n712 VDPWR.n711 0.376971
R3336 VDPWR.n843 VDPWR.n667 0.376971
R3337 VDPWR.n810 VDPWR.n743 0.376971
R3338 VDPWR.n805 VDPWR.n745 0.376971
R3339 VDPWR.n764 VDPWR.n763 0.376971
R3340 VDPWR.n688 VDPWR.n680 0.376971
R3341 VDPWR.n691 VDPWR.n679 0.376971
R3342 VDPWR.n833 VDPWR.n665 0.376971
R3343 VDPWR.n751 VDPWR.n744 0.376971
R3344 VDPWR.n757 VDPWR.n756 0.376971
R3345 VDPWR.n503 VDPWR.n502 0.376971
R3346 VDPWR.n509 VDPWR.n471 0.376971
R3347 VDPWR.n499 VDPWR.n482 0.376971
R3348 VDPWR.n492 VDPWR.n469 0.376971
R3349 VDPWR.n551 VDPWR.n550 0.376971
R3350 VDPWR.n557 VDPWR.n519 0.376971
R3351 VDPWR.n547 VDPWR.n530 0.376971
R3352 VDPWR.n540 VDPWR.n517 0.376971
R3353 VDPWR.n456 VDPWR.n330 0.376971
R3354 VDPWR.n414 VDPWR.n413 0.376971
R3355 VDPWR.n87 VDPWR.n4 0.376971
R3356 VDPWR.n12 VDPWR.n11 0.376971
R3357 VDPWR.n67 VDPWR.n66 0.376971
R3358 VDPWR.n32 VDPWR.n31 0.376971
R3359 VDPWR.n40 VDPWR.n39 0.376971
R3360 VDPWR.n224 VDPWR.n184 0.376971
R3361 VDPWR.n110 VDPWR.n94 0.376971
R3362 VDPWR.n319 VDPWR.n98 0.376971
R3363 VDPWR.n226 VDPWR.n181 0.376971
R3364 VDPWR.n642 VDPWR.n566 0.376971
R3365 VDPWR.n646 VDPWR 0.376726
R3366 VDPWR.n809 VDPWR.n808 0.360656
R3367 VDPWR.n844 VDPWR.n666 0.360656
R3368 VDPWR.n621 VDPWR 0.349949
R3369 VDPWR.n623 VDPWR 0.344944
R3370 VDPWR.n648 VDPWR.n562 0.34097
R3371 VDPWR.n653 VDPWR.n652 0.321157
R3372 VDPWR.n440 VDPWR.n439 0.307571
R3373 VDPWR.n393 VDPWR.n389 0.307571
R3374 VDPWR.n196 VDPWR.n194 0.307571
R3375 VDPWR.n305 VDPWR.n304 0.307571
R3376 VDPWR.n300 VDPWR.n299 0.307571
R3377 VDPWR.n234 VDPWR.n169 0.307571
R3378 VDPWR.n601 VDPWR.n600 0.307571
R3379 VDPWR.n645 VDPWR 0.304352
R3380 VDPWR.n625 VDPWR.n624 0.291125
R3381 VDPWR.n623 VDPWR.n622 0.277007
R3382 VDPWR.n409 VDPWR 0.27355
R3383 VDPWR.n624 VDPWR.n621 0.2731
R3384 VDPWR.n327 VDPWR 0.272663
R3385 VDPWR.n96 VDPWR 0.254776
R3386 VDPWR.n93 VDPWR 0.254776
R3387 VDPWR.n513 VDPWR.n512 0.249058
R3388 VDPWR.n463 VDPWR.n462 0.244984
R3389 VDPWR.n328 VDPWR 0.244503
R3390 VDPWR.n410 VDPWR 0.244503
R3391 VDPWR.n464 VDPWR.n463 0.234803
R3392 VDPWR.n561 VDPWR.n560 0.232427
R3393 VDPWR.n65 VDPWR.n0 0.22821
R3394 VDPWR.n515 VDPWR.n2 0.218931
R3395 VDPWR.n516 VDPWR.n468 0.204432
R3396 VDPWR.n65 VDPWR.n64 0.201986
R3397 VDPWR.n655 VDPWR.n465 0.193242
R3398 VDPWR.n512 VDPWR.n1 0.189404
R3399 VDPWR.n450 VDPWR.n449 0.178728
R3400 VDPWR.n399 VDPWR.n398 0.178728
R3401 VDPWR.n191 VDPWR.n190 0.178728
R3402 VDPWR.n283 VDPWR.n279 0.178728
R3403 VDPWR.n290 VDPWR.n132 0.178728
R3404 VDPWR.n240 VDPWR.n239 0.178728
R3405 VDPWR.n608 VDPWR.n576 0.178728
R3406 VDPWR.n664 VDPWR.n663 0.171208
R3407 VDPWR.n662 VDPWR.n3 0.171141
R3408 VDPWR.n661 VDPWR.n660 0.166741
R3409 VDPWR.n664 VDPWR.n2 0.166514
R3410 VDPWR.n710 VDPWR 0.166125
R3411 VDPWR.n806 VDPWR 0.164562
R3412 VDPWR VDPWR.n708 0.164562
R3413 VDPWR.n501 VDPWR 0.164562
R3414 VDPWR.n549 VDPWR 0.164562
R3415 VDPWR.n515 VDPWR.n514 0.163619
R3416 VDPWR.n468 VDPWR.n467 0.162949
R3417 VDPWR.n651 VDPWR.n650 0.153104
R3418 VDPWR.n654 VDPWR.n466 0.1514
R3419 VDPWR VDPWR.n460 0.148
R3420 VDPWR.n321 VDPWR.n320 0.147704
R3421 VDPWR.n225 VDPWR.n182 0.147704
R3422 VDPWR.n320 VDPWR.n97 0.146059
R3423 VDPWR.n225 VDPWR.n183 0.146059
R3424 VDPWR.n457 VDPWR.n456 0.133357
R3425 VDPWR.n413 VDPWR.n412 0.133357
R3426 VDPWR.n320 VDPWR.n94 0.133357
R3427 VDPWR.n320 VDPWR.n319 0.133357
R3428 VDPWR.n226 VDPWR.n225 0.133357
R3429 VDPWR.n225 VDPWR.n224 0.133357
R3430 VDPWR.n643 VDPWR.n642 0.133357
R3431 VDPWR.n96 VDPWR.n95 0.131257
R3432 VDPWR.n659 VDPWR.n92 0.131257
R3433 VDPWR.n658 VDPWR.n93 0.131257
R3434 VDPWR.n323 VDPWR.n322 0.129612
R3435 VDPWR.n649 VDPWR.n91 0.125788
R3436 VDPWR.n622 VDPWR 0.113524
R3437 VDPWR.n643 VDPWR.n565 0.110181
R3438 VDPWR.n762 VDPWR.n761 0.109875
R3439 VDPWR.n807 VDPWR.n806 0.109875
R3440 VDPWR.n710 VDPWR.n709 0.109875
R3441 VDPWR.n708 VDPWR.n681 0.109875
R3442 VDPWR.n510 VDPWR.n470 0.109875
R3443 VDPWR.n501 VDPWR.n500 0.109875
R3444 VDPWR.n558 VDPWR.n518 0.109875
R3445 VDPWR.n549 VDPWR.n548 0.109875
R3446 VDPWR.n644 VDPWR.n643 0.108956
R3447 VDPWR VDPWR.n323 0.100037
R3448 VDPWR.n646 VDPWR.n645 0.0979265
R3449 VDPWR.n450 VDPWR.n341 0.0977152
R3450 VDPWR.n398 VDPWR.n397 0.0977152
R3451 VDPWR.n218 VDPWR.n191 0.0977152
R3452 VDPWR.n279 VDPWR.n108 0.0977152
R3453 VDPWR.n291 VDPWR.n290 0.0977152
R3454 VDPWR.n239 VDPWR.n238 0.0977152
R3455 VDPWR.n636 VDPWR.n576 0.0977152
R3456 VDPWR.n647 VDPWR.n563 0.096701
R3457 VDPWR.n514 VDPWR.n513 0.0952222
R3458 VDPWR.n663 VDPWR.n1 0.0952222
R3459 VDPWR.n561 VDPWR.n467 0.0952222
R3460 VDPWR VDPWR.n63 0.0931573
R3461 VDPWR VDPWR.n37 0.0922832
R3462 VDPWR.n88 VDPWR 0.0922832
R3463 VDPWR.n663 VDPWR.n662 0.0884817
R3464 VDPWR.n622 VDPWR 0.0847634
R3465 VDPWR.n458 VDPWR.n457 0.079844
R3466 VDPWR.n412 VDPWR.n406 0.079844
R3467 VDPWR.n514 VDPWR.n466 0.0789784
R3468 VDPWR.n457 VDPWR.n329 0.0789574
R3469 VDPWR.n412 VDPWR.n411 0.0789574
R3470 VDPWR.n650 VDPWR.n467 0.078882
R3471 VDPWR.n846 VDPWR.n845 0.0780862
R3472 VDPWR.n847 VDPWR.n1 0.0742538
R3473 VDPWR.n651 VDPWR.n465 0.0715417
R3474 VDPWR.n328 VDPWR.n327 0.0709787
R3475 VDPWR.n460 VDPWR.n459 0.0709787
R3476 VDPWR.n408 VDPWR.n407 0.0709787
R3477 VDPWR.n410 VDPWR.n409 0.0700922
R3478 VDPWR VDPWR.n564 0.0630773
R3479 VDPWR.n656 VDPWR.n655 0.0627018
R3480 VDPWR.n463 VDPWR.n3 0.0625
R3481 VDPWR.n37 VDPWR.n36 0.0616888
R3482 VDPWR.n63 VDPWR.n62 0.0616888
R3483 VDPWR.n89 VDPWR.n88 0.0616888
R3484 VDPWR.n655 VDPWR.n654 0.0573333
R3485 VDPWR.n648 VDPWR.n647 0.0572867
R3486 VDPWR.n761 VDPWR 0.0551875
R3487 VDPWR VDPWR.n807 0.0551875
R3488 VDPWR.n709 VDPWR 0.0551875
R3489 VDPWR.n681 VDPWR 0.0551875
R3490 VDPWR VDPWR.n470 0.0551875
R3491 VDPWR.n500 VDPWR 0.0551875
R3492 VDPWR VDPWR.n518 0.0551875
R3493 VDPWR.n548 VDPWR 0.0551875
R3494 VDPWR.n660 VDPWR.n91 0.0549669
R3495 VDPWR.n461 VDPWR 0.0545625
R3496 VDPWR.n808 VDPWR 0.0512812
R3497 VDPWR VDPWR.n666 0.0512812
R3498 VDPWR.n646 VDPWR.n564 0.045162
R3499 VDPWR.n662 VDPWR.n661 0.043125
R3500 VDPWR.n650 VDPWR.n649 0.03925
R3501 VDPWR.n656 VDPWR.n464 0.0388531
R3502 VDPWR.n466 VDPWR.n91 0.0360208
R3503 VDPWR.n409 VDPWR.n326 0.0351875
R3504 VDPWR.n324 VDPWR 0.0334335
R3505 VDPWR.n658 VDPWR.n657 0.0315396
R3506 VDPWR.n38 VDPWR 0.0310944
R3507 VDPWR.n36 VDPWR 0.0310944
R3508 VDPWR.n62 VDPWR 0.0310944
R3509 VDPWR VDPWR.n89 0.0310944
R3510 VDPWR.n408 VDPWR.n90 0.0298951
R3511 VDPWR.n64 VDPWR 0.0289091
R3512 VDPWR.n327 VDPWR 0.0265417
R3513 VDPWR.n462 VDPWR.n325 0.0256039
R3514 VDPWR.n560 VDPWR.n513 0.0160462
R3515 VDPWR.n516 VDPWR.n515 0.0149983
R3516 VDPWR.n95 VDPWR 0.0140031
R3517 VDPWR.n461 VDPWR.n326 0.008
R3518 VDPWR.n95 VDPWR 0.00744444
R3519 VDPWR VDPWR.n847 0.00538077
R3520 VDPWR.n624 VDPWR.n623 0.00440625
R3521 VDPWR.n325 VDPWR 0.00308012
R3522 VDPWR.n845 VDPWR 0.00284375
R3523 VDPWR.n657 VDPWR.n324 0.00113131
R3524 ua[1].n1 ua[1] 9.55241
R3525 ua[1].n0 ua[1] 2.51601
R3526 ua[1].n0 ua[1] 2.11902
R3527 ua[1].n1 ua[1].n0 0.188289
R3528 ua[1] ua[1].n1 0.0879542
R3529 flashADC_3bit_0/comp_p_1/out_left.n1 flashADC_3bit_0/comp_p_1/out_left.t2 145.612
R3530 flashADC_3bit_0/comp_p_1/out_left.n2 flashADC_3bit_0/comp_p_1/out_left.t0 143.417
R3531 flashADC_3bit_0/comp_p_1/out_left.n0 flashADC_3bit_0/comp_p_1/out_left.t1 29.4286
R3532 flashADC_3bit_0/comp_p_1/out_left flashADC_3bit_0/comp_p_1/out_left.n3 11.6041
R3533 flashADC_3bit_0/comp_p_1/out_left.n3 flashADC_3bit_0/comp_p_1/out_left.n2 4.33076
R3534 flashADC_3bit_0/comp_p_1/out_left.n1 flashADC_3bit_0/comp_p_1/out_left.n0 2.12634
R3535 flashADC_3bit_0/comp_p_1/out_left.n2 flashADC_3bit_0/comp_p_1/out_left.n1 2.04428
R3536 flashADC_3bit_0/comp_p_1/out_left.n3 flashADC_3bit_0/comp_p_1/out_left.n0 0.00290385
R3537 uo_out[3].n0 uo_out[3].t1 556.78
R3538 uo_out[3].t1 uo_out[3] 547.24
R3539 uo_out[3] uo_out[3].t0 372.113
R3540 uo_out[3].n0 uo_out[3] 9.54008
R3541 uo_out[3].n3 uo_out[3].n2 4.55415
R3542 uo_out[3].n2 uo_out[3] 4.43618
R3543 uo_out[3].n3 uo_out[3] 3.33965
R3544 uo_out[3].n1 uo_out[3].n0 0.253625
R3545 uo_out[3] uo_out[3] 0.063
R3546 uo_out[3].n2 uo_out[3] 0.0443144
R3547 uo_out[3] uo_out[3].n3 0.0262742
R3548 uo_out[3] uo_out[3] 0.0262732
R3549 uo_out[3].n1 uo_out[3] 0.013
R3550 uo_out[3].n3 uo_out[3] 0.00801031
R3551 uo_out[3] uo_out[3].n1 0.00565464
R3552 ua[0].n20 ua[0].t26 899.324
R3553 ua[0].n38 ua[0].t22 899.324
R3554 ua[0].n31 ua[0].t14 899.324
R3555 ua[0].n25 ua[0].t2 899.324
R3556 ua[0].n2 ua[0].t6 899.324
R3557 ua[0].n7 ua[0].t10 899.324
R3558 ua[0].n13 ua[0].t18 899.324
R3559 ua[0].n21 ua[0].t26 898.659
R3560 ua[0].n39 ua[0].t22 898.659
R3561 ua[0].n32 ua[0].t14 898.659
R3562 ua[0].n26 ua[0].t2 898.659
R3563 ua[0].n3 ua[0].t6 898.659
R3564 ua[0].n8 ua[0].t10 898.659
R3565 ua[0].n14 ua[0].t18 898.659
R3566 ua[0].t23 ua[0].n38 898.442
R3567 ua[0].t3 ua[0].n25 898.442
R3568 ua[0].t7 ua[0].n2 898.442
R3569 ua[0].t19 ua[0].n13 898.442
R3570 ua[0].t27 ua[0].n20 898.442
R3571 ua[0].t15 ua[0].n31 898.442
R3572 ua[0].t11 ua[0].n7 898.442
R3573 ua[0].n21 ua[0].t27 897.754
R3574 ua[0].n39 ua[0].t23 897.754
R3575 ua[0].n32 ua[0].t15 897.754
R3576 ua[0].n26 ua[0].t3 897.754
R3577 ua[0].n3 ua[0].t7 897.754
R3578 ua[0].n8 ua[0].t11 897.754
R3579 ua[0].n14 ua[0].t19 897.754
R3580 ua[0].n18 ua[0].t24 895.625
R3581 ua[0].n36 ua[0].t20 895.625
R3582 ua[0].n29 ua[0].t12 895.625
R3583 ua[0].n23 ua[0].t0 895.625
R3584 ua[0].n0 ua[0].t4 895.625
R3585 ua[0].n5 ua[0].t8 895.625
R3586 ua[0].n11 ua[0].t16 895.625
R3587 ua[0].n18 ua[0].t25 894.172
R3588 ua[0].n36 ua[0].t21 894.172
R3589 ua[0].n29 ua[0].t13 894.172
R3590 ua[0].n23 ua[0].t1 894.172
R3591 ua[0].n0 ua[0].t5 894.172
R3592 ua[0].n5 ua[0].t9 894.172
R3593 ua[0].n11 ua[0].t17 894.172
R3594 ua[0] ua[0] 11.363
R3595 ua[0].n19 ua[0].n18 6.30807
R3596 ua[0].n37 ua[0].n36 6.30807
R3597 ua[0].n30 ua[0].n29 6.30807
R3598 ua[0].n24 ua[0].n23 6.30807
R3599 ua[0].n1 ua[0].n0 6.30807
R3600 ua[0].n6 ua[0].n5 6.30807
R3601 ua[0].n12 ua[0].n11 6.30807
R3602 ua[0].n20 ua[0].n19 5.39021
R3603 ua[0].n38 ua[0].n37 5.39021
R3604 ua[0].n31 ua[0].n30 5.39021
R3605 ua[0].n25 ua[0].n24 5.39021
R3606 ua[0].n2 ua[0].n1 5.39021
R3607 ua[0].n7 ua[0].n6 5.39021
R3608 ua[0].n13 ua[0].n12 5.39021
R3609 ua[0].n22 ua[0].n21 5.38653
R3610 ua[0].n40 ua[0].n39 5.38653
R3611 ua[0].n33 ua[0].n32 5.38653
R3612 ua[0].n27 ua[0].n26 5.38653
R3613 ua[0].n4 ua[0].n3 5.38653
R3614 ua[0].n9 ua[0].n8 5.38653
R3615 ua[0].n15 ua[0].n14 5.38653
R3616 ua[0].n44 ua[0].n43 5.20469
R3617 ua[0].n22 ua[0].n19 5.11108
R3618 ua[0].n40 ua[0].n37 5.11108
R3619 ua[0].n33 ua[0].n30 5.11108
R3620 ua[0].n27 ua[0].n24 5.11108
R3621 ua[0].n4 ua[0].n1 5.11108
R3622 ua[0].n9 ua[0].n6 5.11108
R3623 ua[0].n15 ua[0].n12 5.11108
R3624 ua[0].n35 ua[0].n28 4.57467
R3625 ua[0].n10 ua[0] 4.13219
R3626 ua[0].n35 ua[0].n34 3.68222
R3627 ua[0].n42 ua[0].n41 3.10272
R3628 ua[0].n16 ua[0] 2.68025
R3629 ua[0].n10 ua[0] 2.66582
R3630 ua[0].n43 ua[0].n42 2.43775
R3631 ua[0].n43 ua[0] 1.54614
R3632 ua[0].n17 ua[0].n16 1.35915
R3633 ua[0] ua[0].n22 0.870692
R3634 ua[0] ua[0].n4 0.870692
R3635 ua[0] ua[0].n9 0.870692
R3636 ua[0] ua[0].n15 0.870692
R3637 ua[0].n34 ua[0].n33 0.837038
R3638 ua[0].n41 ua[0].n40 0.726462
R3639 ua[0].n16 ua[0].n10 0.70492
R3640 ua[0].n28 ua[0].n27 0.668769
R3641 ua[0].n42 ua[0].n35 0.533734
R3642 ua[0].n17 ua[0] 0.468179
R3643 ua[0] ua[0].n45 0.332981
R3644 ua[0].n45 ua[0] 0.20608
R3645 ua[0].n41 ua[0] 0.0482941
R3646 ua[0].n44 ua[0].n17 0.0422977
R3647 ua[0].n45 ua[0].n44 0.0422977
R3648 ua[0].n28 ua[0] 0.0391905
R3649 ua[0].n34 ua[0] 0.0341538
R3650 flashADC_3bit_0/comp_p_0/latch_right.n1 flashADC_3bit_0/comp_p_0/latch_right.t3 114.778
R3651 flashADC_3bit_0/comp_p_0/latch_right.n1 flashADC_3bit_0/comp_p_0/latch_right.t2 106.572
R3652 flashADC_3bit_0/comp_p_0/latch_right.n2 flashADC_3bit_0/comp_p_0/latch_right.t0 94.6192
R3653 flashADC_3bit_0/comp_p_0/latch_right.n0 flashADC_3bit_0/comp_p_0/latch_right.t1 22.0141
R3654 flashADC_3bit_0/comp_p_0/latch_right.n2 flashADC_3bit_0/comp_p_0/latch_right.n0 2.37533
R3655 flashADC_3bit_0/comp_p_0/latch_right.n3 flashADC_3bit_0/comp_p_0/latch_right.n1 1.43373
R3656 flashADC_3bit_0/comp_p_0/latch_right.n4 flashADC_3bit_0/comp_p_0/latch_right.n3 1.11841
R3657 flashADC_3bit_0/comp_p_0/latch_right.n3 flashADC_3bit_0/comp_p_0/latch_right.n2 1.06963
R3658 flashADC_3bit_0/comp_p_0/latch_right flashADC_3bit_0/comp_p_0/latch_right.n4 0.608139
R3659 flashADC_3bit_0/comp_p_0/latch_right.n4 flashADC_3bit_0/comp_p_0/latch_right.n0 0.00530769
R3660 flashADC_3bit_0/comp_p_0/out_left.n1 flashADC_3bit_0/comp_p_0/out_left.t2 145.612
R3661 flashADC_3bit_0/comp_p_0/out_left.n2 flashADC_3bit_0/comp_p_0/out_left.t0 143.417
R3662 flashADC_3bit_0/comp_p_0/out_left.n0 flashADC_3bit_0/comp_p_0/out_left.t1 29.4286
R3663 flashADC_3bit_0/comp_p_0/out_left flashADC_3bit_0/comp_p_0/out_left.n3 11.6041
R3664 flashADC_3bit_0/comp_p_0/out_left.n3 flashADC_3bit_0/comp_p_0/out_left.n2 4.33076
R3665 flashADC_3bit_0/comp_p_0/out_left.n1 flashADC_3bit_0/comp_p_0/out_left.n0 2.12634
R3666 flashADC_3bit_0/comp_p_0/out_left.n2 flashADC_3bit_0/comp_p_0/out_left.n1 2.04428
R3667 flashADC_3bit_0/comp_p_0/out_left.n3 flashADC_3bit_0/comp_p_0/out_left.n0 0.00290385
R3668 uo_out[4].n0 uo_out[4].t1 556.78
R3669 uo_out[4].t1 uo_out[4] 547.24
R3670 uo_out[4] uo_out[4].t0 372.113
R3671 uo_out[4].n1 uo_out[4] 20.4931
R3672 uo_out[4].n0 uo_out[4] 9.54008
R3673 uo_out[4].n2 uo_out[4] 4.35598
R3674 uo_out[4].n2 uo_out[4].n1 3.45922
R3675 uo_out[4].n1 uo_out[4] 1.38807
R3676 uo_out[4] uo_out[4].n0 0.266125
R3677 uo_out[4] uo_out[4] 0.063
R3678 uo_out[4] uo_out[4].n2 0.0217258
R3679 uo_out[4].n2 uo_out[4] 0.00887356
R3680 flashADC_3bit_0/comp_p_2/latch_left.n0 flashADC_3bit_0/comp_p_2/latch_left.t3 114.778
R3681 flashADC_3bit_0/comp_p_2/latch_left.n0 flashADC_3bit_0/comp_p_2/latch_left.t2 106.572
R3682 flashADC_3bit_0/comp_p_2/latch_left.n1 flashADC_3bit_0/comp_p_2/latch_left.t0 95.1712
R3683 flashADC_3bit_0/comp_p_2/latch_left.n2 flashADC_3bit_0/comp_p_2/latch_left.t1 22.0141
R3684 flashADC_3bit_0/comp_p_2/latch_left.n1 flashADC_3bit_0/comp_p_2/latch_left.n0 1.72733
R3685 flashADC_3bit_0/comp_p_2/latch_left flashADC_3bit_0/comp_p_2/latch_left.n2 0.717514
R3686 flashADC_3bit_0/comp_p_2/latch_left.n2 flashADC_3bit_0/comp_p_2/latch_left.n1 0.599169
R3687 uo_out[5].n0 uo_out[5].t1 556.78
R3688 uo_out[5].t1 uo_out[5] 547.24
R3689 uo_out[5] uo_out[5].t0 372.113
R3690 uo_out[5].n2 uo_out[5] 18.5756
R3691 uo_out[5].n0 uo_out[5] 9.54008
R3692 uo_out[5].n3 uo_out[5] 5.91776
R3693 uo_out[5].n2 uo_out[5] 1.06075
R3694 uo_out[5].n3 uo_out[5].n2 0.928508
R3695 uo_out[5].n1 uo_out[5].n0 0.25675
R3696 uo_out[5] uo_out[5].n3 0.0929839
R3697 uo_out[5] uo_out[5] 0.063
R3698 uo_out[5] uo_out[5] 0.0329675
R3699 uo_out[5].n3 uo_out[5] 0.0124426
R3700 uo_out[5].n1 uo_out[5] 0.009875
R3701 uo_out[5] uo_out[5].n1 0.00537013
R3702 uo_out[6].n0 uo_out[6].t1 556.78
R3703 uo_out[6].t1 uo_out[6] 547.24
R3704 uo_out[6] uo_out[6].t0 372.113
R3705 uo_out[6].n1 uo_out[6] 10.0074
R3706 uo_out[6].n0 uo_out[6] 9.54008
R3707 uo_out[6].n3 uo_out[6] 7.20627
R3708 uo_out[6].n2 uo_out[6].n1 1.978
R3709 uo_out[6].n1 uo_out[6] 0.589103
R3710 uo_out[6] uo_out[6].n0 0.266125
R3711 uo_out[6] uo_out[6].n3 0.0975323
R3712 uo_out[6] uo_out[6] 0.063
R3713 uo_out[6].n3 uo_out[6].n2 0.0223063
R3714 uo_out[6].n2 uo_out[6] 0.00579279
R3715 flashADC_3bit_0/comp_p_4/latch_left.n0 flashADC_3bit_0/comp_p_4/latch_left.t3 114.778
R3716 flashADC_3bit_0/comp_p_4/latch_left.n0 flashADC_3bit_0/comp_p_4/latch_left.t2 106.572
R3717 flashADC_3bit_0/comp_p_4/latch_left.n1 flashADC_3bit_0/comp_p_4/latch_left.t0 95.1712
R3718 flashADC_3bit_0/comp_p_4/latch_left.n2 flashADC_3bit_0/comp_p_4/latch_left.t1 22.0141
R3719 flashADC_3bit_0/comp_p_4/latch_left.n1 flashADC_3bit_0/comp_p_4/latch_left.n0 1.72733
R3720 flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/comp_p_4/latch_left.n2 0.717514
R3721 flashADC_3bit_0/comp_p_4/latch_left.n2 flashADC_3bit_0/comp_p_4/latch_left.n1 0.599169
R3722 uo_out[7].n0 uo_out[7].t1 556.78
R3723 uo_out[7].t1 uo_out[7] 547.24
R3724 uo_out[7] uo_out[7].t0 372.113
R3725 uo_out[7].n1 uo_out[7] 24.2927
R3726 uo_out[7].n0 uo_out[7] 9.54008
R3727 uo_out[7].n2 uo_out[7] 8.84384
R3728 uo_out[7].n1 uo_out[7] 1.81119
R3729 uo_out[7].n2 uo_out[7].n1 1.17633
R3730 uo_out[7] uo_out[7].n0 0.266125
R3731 uo_out[7] uo_out[7] 0.063
R3732 uo_out[7].n2 uo_out[7] 0.0115379
R3733 uo_out[7] uo_out[7].n2 0.00656452
R3734 flashADC_3bit_0/comp_p_5/out_left.n1 flashADC_3bit_0/comp_p_5/out_left.t2 145.612
R3735 flashADC_3bit_0/comp_p_5/out_left.n2 flashADC_3bit_0/comp_p_5/out_left.t0 143.417
R3736 flashADC_3bit_0/comp_p_5/out_left.n0 flashADC_3bit_0/comp_p_5/out_left.t1 29.4286
R3737 flashADC_3bit_0/comp_p_5/out_left flashADC_3bit_0/comp_p_5/out_left.n3 11.6041
R3738 flashADC_3bit_0/comp_p_5/out_left.n3 flashADC_3bit_0/comp_p_5/out_left.n2 4.33076
R3739 flashADC_3bit_0/comp_p_5/out_left.n1 flashADC_3bit_0/comp_p_5/out_left.n0 2.12634
R3740 flashADC_3bit_0/comp_p_5/out_left.n2 flashADC_3bit_0/comp_p_5/out_left.n1 2.04428
R3741 flashADC_3bit_0/comp_p_5/out_left.n3 flashADC_3bit_0/comp_p_5/out_left.n0 0.00290385
R3742 uio_out[0].n0 uio_out[0].t1 556.78
R3743 uio_out[0].t1 uio_out[0] 547.24
R3744 uio_out[0] uio_out[0].t0 372.113
R3745 uio_out[0].n2 uio_out[0] 9.82897
R3746 uio_out[0].n0 uio_out[0] 9.54008
R3747 uio_out[0].n2 uio_out[0].n1 3.01518
R3748 uio_out[0].n1 uio_out[0] 2.80934
R3749 uio_out[0].n1 uio_out[0] 0.322375
R3750 uio_out[0] uio_out[0].n0 0.266125
R3751 uio_out[0] uio_out[0] 0.063
R3752 uio_out[0] uio_out[0].n2 0.0213143
R3753 flashADC_3bit_0/comp_p_6/latch_left.n0 flashADC_3bit_0/comp_p_6/latch_left.t3 114.778
R3754 flashADC_3bit_0/comp_p_6/latch_left.n0 flashADC_3bit_0/comp_p_6/latch_left.t2 106.572
R3755 flashADC_3bit_0/comp_p_6/latch_left.n1 flashADC_3bit_0/comp_p_6/latch_left.t0 95.1712
R3756 flashADC_3bit_0/comp_p_6/latch_left.n2 flashADC_3bit_0/comp_p_6/latch_left.t1 22.0141
R3757 flashADC_3bit_0/comp_p_6/latch_left.n1 flashADC_3bit_0/comp_p_6/latch_left.n0 1.72733
R3758 flashADC_3bit_0/comp_p_6/latch_left flashADC_3bit_0/comp_p_6/latch_left.n2 0.717514
R3759 flashADC_3bit_0/comp_p_6/latch_left.n2 flashADC_3bit_0/comp_p_6/latch_left.n1 0.599169
R3760 uio_out[1].n0 uio_out[1].t1 556.78
R3761 uio_out[1].t1 uio_out[1] 547.24
R3762 uio_out[1] uio_out[1].t0 372.113
R3763 uio_out[1].n1 uio_out[1] 11.4942
R3764 uio_out[1].n2 uio_out[1] 11.3634
R3765 uio_out[1].n0 uio_out[1] 9.54008
R3766 uio_out[1].n2 uio_out[1].n1 3.83483
R3767 uio_out[1].n1 uio_out[1] 1.33473
R3768 uio_out[1] uio_out[1].n0 0.266125
R3769 uio_out[1] uio_out[1] 0.063
R3770 uio_out[1] uio_out[1].n2 0.0550806
R3771 uio_out[1].n2 uio_out[1] 0.0207361
R3772 uo_out[0].n0 uo_out[0] 8.08738
R3773 uo_out[0].n0 uo_out[0] 5.30089
R3774 uo_out[0].n0 uo_out[0] 2.61734
R3775 uo_out[0] uo_out[0].n0 0.03175
R3776 uo_out[1] uo_out[1].n0 9.33705
R3777 uo_out[1].n0 uo_out[1] 5.30089
R3778 uo_out[1].n0 uo_out[1] 2.61734
R3779 uo_out[1].n0 uo_out[1] 0.03175
R3780 uo_out[2] uo_out[2].n0 10.6421
R3781 uo_out[2].n0 uo_out[2] 5.30089
R3782 uo_out[2].n0 uo_out[2] 2.61734
R3783 uo_out[2].n0 uo_out[2] 0.03175
C0 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_3/vinn -0.01472f
C1 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out 1.04758f
C2 VDPWR flashADC_3bit_0/comp_p_1/latch_right 0.22258f
C3 flashADC_3bit_0/comp_p_4/vinn ua[0] -0
C4 VDPWR flashADC_3bit_0/comp_p_2/vinn 0.04885f
C5 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin -0
C6 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out 0.00956f
C7 uo_out[2] uo_out[3] 0.09111f
C8 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B VDPWR 0.21063f
C9 uo_out[4] flashADC_3bit_0/comp_p_3/vinn -0
C10 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_4/tail -0.04111f
C11 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in -0
C12 uo_out[5] flashADC_3bit_0/comp_p_3/vinn -0.00952f
C13 flashADC_3bit_0/comp_p_5/out_left VDPWR 0.47743f
C14 uo_out[4] uo_out[6] 0
C15 uio_oe[3] VDPWR 0
C16 uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin 0.00138f
C17 uio_out[5] VDPWR 0
C18 flashADC_3bit_0/comp_p_1/tail uio_out[1] 0
C19 uio_out[0] uo_out[7] 0.99679f
C20 flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_3/vinn -0.01138f
C21 flashADC_3bit_0/comp_p_0/vinn VDPWR 1.85762f
C22 flashADC_3bit_0/comp_p_4/out_left flashADC_3bit_0/comp_p_5/vinn -0.00479f
C23 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin -0
C24 uo_out[5] uo_out[6] 0.83351f
C25 flashADC_3bit_0/comp_p_1/vinn VDPWR 1.17123f
C26 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin 0
C27 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A 0.00574f
C28 VDPWR flashADC_3bit_0/comp_p_1/tail 0.02796f
C29 uio_in[2] uio_in[1] 0.03102f
C30 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0.01579f
C31 VDPWR flashADC_3bit_0/comp_p_5/latch_left 0.38506f
C32 uo_out[5] uio_out[1] 0
C33 ua[0] flashADC_3bit_0/comp_p_5/vinn -0.04026f
C34 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin VDPWR 0.01661f
C35 uio_oe[4] uio_oe[3] 0.03102f
C36 uio_oe[0] uio_oe[1] 0.03102f
C37 uio_out[6] uio_out[5] 0.03102f
C38 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_0/latch_right -0.0159f
C39 uo_out[4] VDPWR 0.65166f
C40 uo_out[3] uo_out[0] 0
C41 flashADC_3bit_0/comp_p_5/vinn uo_out[7] -0.01219f
C42 VDPWR uo_out[5] 1.25716f
C43 uio_oe[2] VDPWR 0
C44 VDPWR flashADC_3bit_0/comp_p_2/tail 0.00107f
C45 VDPWR flashADC_3bit_0/comp_p_3/tail 0.03261f
C46 VDPWR flashADC_3bit_0/comp_p_5/tail 0.78378f
C47 rst_n clk 0.03102f
C48 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin VDPWR 0.0016f
C49 VDPWR flashADC_3bit_0/comp_p_6/latch_left 0.42219f
C50 ua[0] flashADC_3bit_0/comp_p_3/vinn -0.02041f
C51 flashADC_3bit_0/comp_p_0/latch_left VDPWR 0.16971f
C52 flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 VDPWR 0.03356f
C53 flashADC_3bit_0/comp_p_6/out_left VDPWR 0.26382f
C54 VDPWR flashADC_3bit_0/comp_p_4/tail 0.66705f
C55 ua[1] ua[0] 4.5498f
C56 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0.0018f
C57 flashADC_3bit_0/vbias_generation_0/bias_n VDPWR 0.10568f
C58 uio_oe[7] VDPWR 0
C59 flashADC_3bit_0/comp_p_4/out_left VDPWR 0.36618f
C60 uio_oe[1] VDPWR 0
C61 uo_out[7] uo_out[6] 0.83703f
C62 uio_in[4] uo_out[1] 0.01025f
C63 flashADC_3bit_0/comp_p_0/vinn flashADC_3bit_0/comp_p_1/vinn -0.00292f
C64 uio_in[6] uo_out[0] 0.01741f
C65 ua[1] ua[7] 0.01625f
C66 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out uo_out[1] 0
C67 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3] 0
C68 uio_in[1] uio_in[0] 0.03102f
C69 uo_out[2] uo_out[6] 0
C70 uio_out[1] uo_out[7] 0
C71 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in uo_out[1] 0.00492f
C72 flashADC_3bit_0/comp_p_1/out_left uo_out[7] 0
C73 VDPWR ua[0] 6.62902f
C74 uio_out[0] uo_out[3] 0.00111f
C75 VDPWR uo_out[1] 0.017f
C76 uio_out[0] flashADC_3bit_0/comp_p_6/vbias_p 0
C77 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VDPWR 0.87869f
C78 uio_oe[3] uio_oe[2] 0.03102f
C79 uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out 0
C80 flashADC_3bit_0/comp_p_1/vinn uo_out[4] -0.01018f
C81 flashADC_3bit_0/comp_p_2/latch_left flashADC_3bit_0/comp_p_3/vinn -0.00981f
C82 VDPWR uo_out[7] 1.68424f
C83 flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/comp_p_3/vinn -0.00404f
C84 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in uo_out[1] 0.00251f
C85 flashADC_3bit_0/comp_p_1/vinn uo_out[5] -0.0012f
C86 uio_oe[6] VDPWR 0
C87 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G VDPWR 0.0124f
C88 uio_in[5] uo_out[0] 0.01741f
C89 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out VDPWR 1.28865f
C90 ua[1] ua[6] 0.01737f
C91 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in uo_out[2] 0
C92 uo_out[5] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C93 VDPWR uo_out[2] 0.08501f
C94 flashADC_3bit_0/comp_p_3/out_left VDPWR 0.18333f
C95 flashADC_3bit_0/comp_p_0/latch_left flashADC_3bit_0/comp_p_1/vinn -0.01177f
C96 uo_out[4] uo_out[5] 0.69387f
C97 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in uo_out[2] 0
C98 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_6/vbias_p -0.0296f
C99 flashADC_3bit_0/comp_p_6/vinn flashADC_3bit_0/comp_p_5/vinn -0.01917f
C100 uo_out[2] uio_in[3] 0.00766f
C101 ui_in[6] ui_in[5] 0.03102f
C102 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B uo_out[1] 0
C103 flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_5/vinn -0.04257f
C104 flashADC_3bit_0/comp_p_2/latch_left VDPWR 0.20391f
C105 uio_oe[5] VDPWR 0
C106 VDPWR flashADC_3bit_0/comp_p_2/out_left 0.14457f
C107 ui_in[7] ui_in[6] 0.03102f
C108 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out uo_out[0] 0
C109 flashADC_3bit_0/comp_p_3/latch_left VDPWR 0.27789f
C110 flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_3/vinn -0.02616f
C111 flashADC_3bit_0/comp_p_6/tail VDPWR 0.00165f
C112 flashADC_3bit_0/comp_p_0/vinn ua[0] -0
C113 uio_in[0] ui_in[7] 0.03102f
C114 flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/comp_p_5/vinn -0.02278f
C115 clk ena 0.03102f
C116 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B uo_out[2] 0
C117 flashADC_3bit_0/comp_p_1/vinn ua[0] -0.00683f
C118 uo_out[3] uo_out[6] 0
C119 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin uo_out[1] 0.00282f
C120 VDPWR uo_out[0] 0.10165f
C121 uio_oe[4] uio_oe[5] 0.03102f
C122 uio_oe[2] uio_oe[1] 0.03102f
C123 uio_in[2] uio_in[3] 0.03102f
C124 flashADC_3bit_0/comp_p_6/vinn ua[1] 0.19732f
C125 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in uo_out[0] 0.00561f
C126 ui_in[2] ui_in[1] 0.03102f
C127 uio_in[6] uio_in[5] 0.03102f
C128 VDPWR flashADC_3bit_0/comp_p_0/tail 0
C129 uio_out[1] uo_out[3] 0.00552f
C130 flashADC_3bit_0/comp_p_4/latch_right flashADC_3bit_0/comp_p_5/vinn -0.02778f
C131 uio_in[7] uo_out[0] 0.04843f
C132 uio_out[1] flashADC_3bit_0/comp_p_6/vbias_p 0.00692f
C133 uio_out[4] uio_out[3] 0.03102f
C134 ua[5] ua[1] 0.01737f
C135 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin uo_out[2] 0
C136 uo_out[4] uo_out[7] 0
C137 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A uo_out[2] 0
C138 VDPWR uo_out[3] 0.20792f
C139 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_3/vinn -0.01316f
C140 VDPWR flashADC_3bit_0/comp_p_6/vbias_p 5.47005f
C141 uo_out[5] uo_out[7] 0.00111f
C142 flashADC_3bit_0/comp_p_6/vinn VDPWR 0.75805f
C143 uio_out[0] uo_out[6] 0
C144 ui_in[5] ui_in[4] 0.03102f
C145 uo_out[4] uo_out[2] 0
C146 flashADC_3bit_0/comp_p_4/vinn VDPWR 0.57174f
C147 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin 0.00218f
C148 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_2/latch_left -0.00559f
C149 uo_out[5] uo_out[2] 0
C150 flashADC_3bit_0/comp_p_5/latch_right VDPWR 0.3836f
C151 uio_out[0] uio_out[1] 0.94888f
C152 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_3/vinn -0.02012f
C153 uio_out[0] flashADC_3bit_0/comp_p_1/out_left 0
C154 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0.01085f
C155 ua[4] ua[1] 0.01737f
C156 ui_in[2] ui_in[3] 0.03102f
C157 flashADC_3bit_0/comp_p_4/latch_left VDPWR 0.25376f
C158 uio_out[0] VDPWR 1.07221f
C159 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out VDPWR 0.12659f
C160 flashADC_3bit_0/comp_p_2/latch_right VDPWR 0.23507f
C161 VDPWR uio_in[6] 0
C162 VDPWR uio_out[4] 0
C163 uio_oe[7] uio_oe[6] 0.03102f
C164 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A uo_out[0] 0
C165 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin uo_out[1] 0.00143f
C166 ui_in[1] ui_in[0] 0.03102f
C167 uio_in[5] uio_in[4] 0.03102f
C168 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/m1_n100_n100# VDPWR 0.00545f
C169 flashADC_3bit_0/comp_p_4/latch_right VDPWR 0.29499f
C170 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 uo_out[1] 0
C171 uio_in[7] uio_in[6] 0.03102f
C172 ua[0] uo_out[7] -0
C173 uio_out[3] uio_out[2] 0.03102f
C174 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G 0.10354f
C175 ua[3] ua[1] 0.01737f
C176 VDPWR flashADC_3bit_0/comp_p_5/vinn 3.18346f
C177 flashADC_3bit_0/comp_p_0/out_left VDPWR 0.12984f
C178 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_6/vbias_p -0.00683f
C179 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin uo_out[2] 0
C180 VDPWR uio_in[5] 0
C181 uo_out[2] uo_out[1] 2.07257f
C182 VDPWR uio_out[3] 0
C183 uio_oe[0] uio_out[7] 0.03102f
C184 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 uo_out[2] 0.00393f
C185 ui_in[4] ui_in[3] 0.03102f
C186 uo_out[2] uo_out[7] 0
C187 uo_out[1] flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G 0
C188 uo_out[4] uo_out[3] 0.31058f
C189 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 VDPWR 0.0044f
C190 uio_oe[0] VDPWR 0
C191 VDPWR flashADC_3bit_0/comp_p_3/vinn 1.60219f
C192 uo_out[5] uo_out[3] 0
C193 uio_out[1] uo_out[6] 0
C194 ua[2] ua[1] 0.01737f
C195 uio_out[1] uio_out[2] 0.03102f
C196 VDPWR uo_out[6] 0.59661f
C197 uio_out[5] uio_out[4] 0.03102f
C198 ua[1] VDPWR 0.29111f
C199 VDPWR flashADC_3bit_0/comp_p_6/latch_right 0.39269f
C200 uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G 0
C201 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_1/vinn -0.00771f
C202 flashADC_3bit_0/comp_p_1/out_left uio_out[1] 0.03149f
C203 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out 0.45869f
C204 VDPWR uio_out[2] 0
C205 uio_oe[6] uio_oe[5] 0.03102f
C206 VDPWR uio_out[1] 2.03753f
C207 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G VDPWR 0.01001f
C208 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin uo_out[0] 0.00613f
C209 uio_out[7] VDPWR 0
C210 VDPWR flashADC_3bit_0/comp_p_1/out_left 0.15235f
C211 ui_in[0] rst_n 0.03102f
C212 VDPWR flashADC_3bit_0/comp_p_1/latch_left 0.23151f
C213 uio_in[4] uio_in[3] 0.03102f
C214 flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_3/vinn -0.01451f
C215 uo_out[0] uo_out[1] 1.70165f
C216 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VDPWR 0.02718f
C217 VDPWR flashADC_3bit_0/comp_p_3/latch_right 0.26506f
C218 uio_out[0] uo_out[5] 0
C219 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in 0
C220 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_0/out_left -0.00559f
C221 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in VDPWR 0.01474f
C222 VDPWR uio_in[7] 0
C223 uio_out[7] uio_out[6] 0.03102f
C224 uo_out[2] uo_out[0] 0.0867f
C225 VDPWR flashADC_3bit_0/comp_p_0/latch_right 0.19561f
C226 uo_out[3] uo_out[1] 0
C227 flashADC_3bit_0/comp_p_0/vinn flashADC_3bit_0/comp_p_3/vinn -0.03853f
C228 flashADC_3bit_0/comp_p_6/vinn ua[0] 0
C229 uo_out[3] uo_out[7] 0
C230 uio_oe[4] VDPWR 0
C231 uio_out[6] VDPWR 0
C232 ua[2] VGND 0.12712f
C233 ua[3] VGND 0.12712f
C234 ua[4] VGND 0.12712f
C235 ua[5] VGND 0.12712f
C236 ua[6] VGND 0.12712f
C237 ua[7] VGND 0.12842f
C238 ena VGND 0.07038f
C239 clk VGND 0.04288f
C240 rst_n VGND 0.04288f
C241 ui_in[0] VGND 0.04288f
C242 ui_in[1] VGND 0.04288f
C243 ui_in[2] VGND 0.04288f
C244 ui_in[3] VGND 0.04288f
C245 ui_in[4] VGND 0.04288f
C246 ui_in[5] VGND 0.04288f
C247 ui_in[6] VGND 0.04288f
C248 ui_in[7] VGND 0.04288f
C249 uio_in[0] VGND 0.04288f
C250 uio_in[1] VGND 0.04288f
C251 uio_in[2] VGND 0.04288f
C252 uio_in[3] VGND 0.03541f
C253 uio_in[4] VGND 0.03434f
C254 uio_in[5] VGND 0.0331f
C255 uio_in[6] VGND 0.0331f
C256 uio_in[7] VGND 0.0331f
C257 uio_out[2] VGND 0.04167f
C258 uio_out[3] VGND 0.04167f
C259 uio_out[4] VGND 0.04167f
C260 uio_out[5] VGND 0.04167f
C261 uio_out[6] VGND 0.04167f
C262 uio_out[7] VGND 0.04167f
C263 uio_oe[0] VGND 0.04176f
C264 uio_oe[1] VGND 0.04176f
C265 uio_oe[2] VGND 0.04167f
C266 uio_oe[3] VGND 0.04167f
C267 uio_oe[4] VGND 0.04167f
C268 uio_oe[5] VGND 0.04167f
C269 uio_oe[6] VGND 0.04167f
C270 uio_oe[7] VGND 0.06927f
C271 uo_out[2].n0 VGND 0.80677f
C272 uo_out[1].n0 VGND 0.8648f
C273 uio_out[1].t1 VGND 0.09868f
C274 uio_out[1].t0 VGND 0.09363f
C275 uio_out[1].n0 VGND 0.27936f
C276 uio_out[1].n1 VGND 2.99315f
C277 uio_out[1].n2 VGND 4.58739f
C278 flashADC_3bit_0/comp_p_6/latch_left.t0 VGND 1.2884f
C279 flashADC_3bit_0/comp_p_6/latch_left.t3 VGND 1.61523f
C280 flashADC_3bit_0/comp_p_6/latch_left.t2 VGND 1.50002f
C281 flashADC_3bit_0/comp_p_6/latch_left.n0 VGND 2.85187f
C282 flashADC_3bit_0/comp_p_6/latch_left.n1 VGND 1.83029f
C283 flashADC_3bit_0/comp_p_6/latch_left.t1 VGND 0.38521f
C284 flashADC_3bit_0/comp_p_6/latch_left.n2 VGND 1.64625f
C285 uio_out[0].t0 VGND 0.12278f
C286 uio_out[0].t1 VGND 0.1294f
C287 uio_out[0].n0 VGND 0.36633f
C288 uio_out[0].n1 VGND 0.92016f
C289 uio_out[0].n2 VGND 5.10634f
C290 flashADC_3bit_0/comp_p_5/out_left.t1 VGND 0.38277f
C291 flashADC_3bit_0/comp_p_5/out_left.n0 VGND 0.38383f
C292 flashADC_3bit_0/comp_p_5/out_left.t2 VGND 1.01962f
C293 flashADC_3bit_0/comp_p_5/out_left.n1 VGND 1.84849f
C294 flashADC_3bit_0/comp_p_5/out_left.t0 VGND 1.01131f
C295 flashADC_3bit_0/comp_p_5/out_left.n2 VGND 0.33514f
C296 flashADC_3bit_0/comp_p_5/out_left.n3 VGND 1.32622f
C297 uo_out[7].t1 VGND 0.07979f
C298 uo_out[7].t0 VGND 0.07571f
C299 uo_out[7].n0 VGND 0.22588f
C300 uo_out[7].n1 VGND 4.90541f
C301 uo_out[7].n2 VGND 2.61036f
C302 flashADC_3bit_0/comp_p_4/latch_left.t0 VGND 1.01079f
C303 flashADC_3bit_0/comp_p_4/latch_left.t3 VGND 1.2672f
C304 flashADC_3bit_0/comp_p_4/latch_left.t2 VGND 1.17681f
C305 flashADC_3bit_0/comp_p_4/latch_left.n0 VGND 2.23738f
C306 flashADC_3bit_0/comp_p_4/latch_left.n1 VGND 1.43592f
C307 flashADC_3bit_0/comp_p_4/latch_left.t1 VGND 0.30221f
C308 flashADC_3bit_0/comp_p_4/latch_left.n2 VGND 1.29154f
C309 uo_out[6].t0 VGND 0.10769f
C310 uo_out[6].t1 VGND 0.11349f
C311 uo_out[6].n0 VGND 0.3213f
C312 uo_out[6].n1 VGND 2.49197f
C313 uo_out[6].n2 VGND 0.38414f
C314 uo_out[6].n3 VGND 2.88453f
C315 uo_out[5].t1 VGND 0.09276f
C316 uo_out[5].t0 VGND 0.08802f
C317 uo_out[5].n0 VGND 0.26072f
C318 uo_out[5].n1 VGND 0.05704f
C319 uo_out[5].n2 VGND 3.66875f
C320 uo_out[5].n3 VGND 2.20196f
C321 flashADC_3bit_0/comp_p_2/latch_left.t0 VGND 1.01079f
C322 flashADC_3bit_0/comp_p_2/latch_left.t3 VGND 1.2672f
C323 flashADC_3bit_0/comp_p_2/latch_left.t2 VGND 1.17681f
C324 flashADC_3bit_0/comp_p_2/latch_left.n0 VGND 2.23738f
C325 flashADC_3bit_0/comp_p_2/latch_left.n1 VGND 1.43592f
C326 flashADC_3bit_0/comp_p_2/latch_left.t1 VGND 0.30221f
C327 flashADC_3bit_0/comp_p_2/latch_left.n2 VGND 1.29154f
C328 uo_out[4].t0 VGND 0.06216f
C329 uo_out[4].t1 VGND 0.06551f
C330 uo_out[4].n0 VGND 0.18546f
C331 uo_out[4].n1 VGND 2.98325f
C332 uo_out[4].n2 VGND 1.11497f
C333 flashADC_3bit_0/comp_p_0/out_left.t1 VGND 0.27049f
C334 flashADC_3bit_0/comp_p_0/out_left.n0 VGND 0.27124f
C335 flashADC_3bit_0/comp_p_0/out_left.t2 VGND 0.72053f
C336 flashADC_3bit_0/comp_p_0/out_left.n1 VGND 1.30626f
C337 flashADC_3bit_0/comp_p_0/out_left.t0 VGND 0.71466f
C338 flashADC_3bit_0/comp_p_0/out_left.n2 VGND 0.23684f
C339 flashADC_3bit_0/comp_p_0/out_left.n3 VGND 0.9372f
C340 flashADC_3bit_0/comp_p_0/latch_right.t1 VGND 0.38673f
C341 flashADC_3bit_0/comp_p_0/latch_right.n0 VGND 0.76282f
C342 flashADC_3bit_0/comp_p_0/latch_right.t3 VGND 1.62161f
C343 flashADC_3bit_0/comp_p_0/latch_right.t2 VGND 1.50595f
C344 flashADC_3bit_0/comp_p_0/latch_right.n1 VGND 2.57607f
C345 flashADC_3bit_0/comp_p_0/latch_right.t0 VGND 1.2913f
C346 flashADC_3bit_0/comp_p_0/latch_right.n2 VGND 0.3778f
C347 flashADC_3bit_0/comp_p_0/latch_right.n3 VGND 1.70107f
C348 flashADC_3bit_0/comp_p_0/latch_right.n4 VGND 0.23787f
C349 ua[0].t4 VGND 0.35773f
C350 ua[0].t5 VGND 0.35749f
C351 ua[0].n0 VGND 0.48033f
C352 ua[0].n1 VGND 0.37605f
C353 ua[0].t6 VGND 0.26587f
C354 ua[0].n2 VGND 0.43251f
C355 ua[0].t7 VGND 0.26553f
C356 ua[0].n3 VGND 0.42523f
C357 ua[0].n4 VGND 0.20155f
C358 ua[0].t8 VGND 0.35773f
C359 ua[0].t9 VGND 0.35749f
C360 ua[0].n5 VGND 0.48033f
C361 ua[0].n6 VGND 0.37605f
C362 ua[0].t10 VGND 0.26587f
C363 ua[0].n7 VGND 0.43251f
C364 ua[0].t11 VGND 0.26553f
C365 ua[0].n8 VGND 0.42523f
C366 ua[0].n9 VGND 0.20155f
C367 ua[0].n10 VGND 2.95964f
C368 ua[0].t16 VGND 0.35773f
C369 ua[0].t17 VGND 0.35749f
C370 ua[0].n11 VGND 0.48033f
C371 ua[0].n12 VGND 0.37605f
C372 ua[0].t18 VGND 0.26587f
C373 ua[0].n13 VGND 0.43251f
C374 ua[0].t19 VGND 0.26553f
C375 ua[0].n14 VGND 0.42523f
C376 ua[0].n15 VGND 0.20155f
C377 ua[0].n16 VGND 1.90625f
C378 ua[0].n17 VGND 1.60944f
C379 ua[0].t24 VGND 0.35773f
C380 ua[0].t25 VGND 0.35749f
C381 ua[0].n18 VGND 0.48033f
C382 ua[0].n19 VGND 0.37605f
C383 ua[0].t26 VGND 0.26587f
C384 ua[0].n20 VGND 0.43251f
C385 ua[0].t27 VGND 0.26553f
C386 ua[0].n21 VGND 0.42523f
C387 ua[0].n22 VGND 0.20155f
C388 ua[0].t0 VGND 0.35773f
C389 ua[0].t1 VGND 0.35749f
C390 ua[0].n23 VGND 0.48033f
C391 ua[0].n24 VGND 0.37605f
C392 ua[0].t2 VGND 0.26587f
C393 ua[0].n25 VGND 0.43251f
C394 ua[0].t3 VGND 0.26553f
C395 ua[0].n26 VGND 0.42523f
C396 ua[0].n27 VGND 0.19504f
C397 ua[0].n28 VGND 0.91535f
C398 ua[0].t12 VGND 0.35773f
C399 ua[0].t13 VGND 0.35749f
C400 ua[0].n29 VGND 0.48033f
C401 ua[0].n30 VGND 0.37605f
C402 ua[0].t14 VGND 0.26587f
C403 ua[0].n31 VGND 0.43251f
C404 ua[0].t15 VGND 0.26553f
C405 ua[0].n32 VGND 0.42523f
C406 ua[0].n33 VGND 0.20046f
C407 ua[0].n34 VGND 0.20563f
C408 ua[0].n35 VGND 3.05495f
C409 ua[0].t20 VGND 0.35773f
C410 ua[0].t21 VGND 0.35749f
C411 ua[0].n36 VGND 0.48033f
C412 ua[0].n37 VGND 0.37605f
C413 ua[0].t22 VGND 0.26587f
C414 ua[0].n38 VGND 0.43251f
C415 ua[0].t23 VGND 0.26553f
C416 ua[0].n39 VGND 0.42523f
C417 ua[0].n40 VGND 0.1969f
C418 ua[0].n41 VGND 0.26684f
C419 ua[0].n42 VGND 2.37573f
C420 ua[0].n43 VGND 2.18604f
C421 ua[0].n44 VGND 1.16689f
C422 ua[0].n45 VGND 0.81445f
C423 uo_out[3].t1 VGND 0.06421f
C424 uo_out[3].t0 VGND 0.06093f
C425 uo_out[3].n0 VGND 0.18004f
C426 uo_out[3].n1 VGND 0.04119f
C427 uo_out[3].n2 VGND 1.07213f
C428 uo_out[3].n3 VGND 1.08672f
C429 flashADC_3bit_0/comp_p_1/out_left.t1 VGND 0.36236f
C430 flashADC_3bit_0/comp_p_1/out_left.n0 VGND 0.36336f
C431 flashADC_3bit_0/comp_p_1/out_left.t2 VGND 0.96524f
C432 flashADC_3bit_0/comp_p_1/out_left.n1 VGND 1.7499f
C433 flashADC_3bit_0/comp_p_1/out_left.t0 VGND 0.95737f
C434 flashADC_3bit_0/comp_p_1/out_left.n2 VGND 0.31727f
C435 flashADC_3bit_0/comp_p_1/out_left.n3 VGND 1.25549f
C436 ua[1].n0 VGND 0.50626f
C437 ua[1].n1 VGND 2.58175f
C438 VDPWR.n0 VGND 0.44659f
C439 VDPWR.n1 VGND 0.65213f
C440 VDPWR.n2 VGND 1.31109f
C441 VDPWR.n3 VGND 13.2158f
C442 VDPWR.n4 VGND 0.0078f
C443 VDPWR.n5 VGND 0.01556f
C444 VDPWR.n6 VGND 0.12519f
C445 VDPWR.n7 VGND 0.01519f
C446 VDPWR.n8 VGND 0.11428f
C447 VDPWR.n9 VGND 0.01556f
C448 VDPWR.n10 VGND 0.01556f
C449 VDPWR.n11 VGND 0.00544f
C450 VDPWR.n12 VGND 0.0078f
C451 VDPWR.n13 VGND 0.11428f
C452 VDPWR.n14 VGND 0.0101f
C453 VDPWR.n15 VGND 0.0101f
C454 VDPWR.n16 VGND 0.0101f
C455 VDPWR.n17 VGND 0.01024f
C456 VDPWR.n18 VGND 0.00976f
C457 VDPWR.n19 VGND 0.00976f
C458 VDPWR.n20 VGND 0.00976f
C459 VDPWR.n21 VGND 0.11428f
C460 VDPWR.n22 VGND 0.11428f
C461 VDPWR.n23 VGND 0.00976f
C462 VDPWR.n24 VGND 0.01024f
C463 VDPWR.n25 VGND 0.00976f
C464 VDPWR.n26 VGND 0.01519f
C465 VDPWR.n27 VGND 0.01519f
C466 VDPWR.n28 VGND 0.11428f
C467 VDPWR.n29 VGND 0.01556f
C468 VDPWR.n30 VGND 0.01556f
C469 VDPWR.n31 VGND 0.00544f
C470 VDPWR.n32 VGND 0.0078f
C471 VDPWR.n33 VGND 0.12519f
C472 VDPWR.n34 VGND 0.01556f
C473 VDPWR.n35 VGND 0.01556f
C474 VDPWR.n36 VGND 0.07271f
C475 VDPWR.n37 VGND 0.0432f
C476 VDPWR.n38 VGND 0.1401f
C477 VDPWR.n39 VGND 0.00765f
C478 VDPWR.n40 VGND 0.0078f
C479 VDPWR.n42 VGND 0.09975f
C480 VDPWR.n43 VGND 0.01519f
C481 VDPWR.n44 VGND 0.01517f
C482 VDPWR.n45 VGND 0.01519f
C483 VDPWR.n46 VGND 0.09475f
C484 VDPWR.n47 VGND 0.09475f
C485 VDPWR.n48 VGND 0.01519f
C486 VDPWR.n49 VGND 0.01519f
C487 VDPWR.n50 VGND 0.01517f
C488 VDPWR.n51 VGND 0.01519f
C489 VDPWR.n52 VGND 0.47664f
C490 VDPWR.n53 VGND 0.47664f
C491 VDPWR.n54 VGND 0.0101f
C492 VDPWR.n55 VGND 0.11428f
C493 VDPWR.n56 VGND 0.0101f
C494 VDPWR.n57 VGND 0.0101f
C495 VDPWR.n58 VGND 0.01024f
C496 VDPWR.n59 VGND 0.01024f
C497 VDPWR.n60 VGND 0.00976f
C498 VDPWR.n61 VGND 0.00974f
C499 VDPWR.n62 VGND 0.07271f
C500 VDPWR.n63 VGND 0.04345f
C501 VDPWR.n64 VGND 0.11484f
C502 VDPWR.n65 VGND 0.1212f
C503 VDPWR.n66 VGND 0.00232f
C504 VDPWR.n67 VGND 0.00233f
C505 VDPWR.n68 VGND 0.00464f
C506 VDPWR.n69 VGND 0.11428f
C507 VDPWR.n70 VGND 0.00464f
C508 VDPWR.n71 VGND 0.00976f
C509 VDPWR.n72 VGND 0.01519f
C510 VDPWR.n73 VGND 0.01519f
C511 VDPWR.n74 VGND 0.09547f
C512 VDPWR.n75 VGND 0.09547f
C513 VDPWR.n76 VGND 0.01519f
C514 VDPWR.n77 VGND 0.01519f
C515 VDPWR.n78 VGND 0.01517f
C516 VDPWR.n79 VGND 0.01519f
C517 VDPWR.n80 VGND 0.09475f
C518 VDPWR.n81 VGND 0.09475f
C519 VDPWR.n82 VGND 0.01519f
C520 VDPWR.n83 VGND 0.01556f
C521 VDPWR.n85 VGND 0.09975f
C522 VDPWR.n86 VGND 0.01517f
C523 VDPWR.n87 VGND 0.00544f
C524 VDPWR.n88 VGND 0.0432f
C525 VDPWR.n89 VGND 0.07271f
C526 VDPWR.n90 VGND 1.12405f
C527 VDPWR.n91 VGND 1.73744f
C528 VDPWR.n92 VGND 0.51583f
C529 VDPWR.n93 VGND 0.36178f
C530 VDPWR.n94 VGND 0.01417f
C531 VDPWR.n95 VGND 0.08035f
C532 VDPWR.n96 VGND 0.36178f
C533 VDPWR.n97 VGND 0.39028f
C534 VDPWR.n98 VGND 0.0175f
C535 VDPWR.n99 VGND 0.21034f
C536 VDPWR.n100 VGND 0.03166f
C537 VDPWR.n101 VGND 0.03579f
C538 VDPWR.n102 VGND 2.23761f
C539 VDPWR.n103 VGND 0.03176f
C540 VDPWR.n104 VGND 0.03176f
C541 VDPWR.n105 VGND 0.40313f
C542 VDPWR.n106 VGND 0.03166f
C543 VDPWR.n107 VGND 0.03579f
C544 VDPWR.n108 VGND 0.11558f
C545 VDPWR.n109 VGND -0.08114f
C546 VDPWR.n110 VGND 0.0175f
C547 VDPWR.n111 VGND 0.03579f
C548 VDPWR.n112 VGND 0.02932f
C549 VDPWR.n113 VGND 0.50278f
C550 VDPWR.n114 VGND 0.03176f
C551 VDPWR.n115 VGND 2.18778f
C552 VDPWR.n116 VGND 0.03176f
C553 VDPWR.n117 VGND 0.10692f
C554 VDPWR.n118 VGND 0.20856f
C555 VDPWR.n119 VGND 0.65798f
C556 VDPWR.n120 VGND 0.04101f
C557 VDPWR.n121 VGND 0.04101f
C558 VDPWR.n122 VGND 2.45276f
C559 VDPWR.n123 VGND 0.04101f
C560 VDPWR.n124 VGND 0.04101f
C561 VDPWR.n125 VGND 0.02932f
C562 VDPWR.n126 VGND 0.03579f
C563 VDPWR.n127 VGND 0.20856f
C564 VDPWR.n128 VGND 0.65798f
C565 VDPWR.n129 VGND 0.10692f
C566 VDPWR.n130 VGND 0.10617f
C567 VDPWR.n131 VGND 0.11454f
C568 VDPWR.n132 VGND 0.37059f
C569 VDPWR.n133 VGND 0.04078f
C570 VDPWR.n134 VGND 0.04093f
C571 VDPWR.n135 VGND 0.67366f
C572 VDPWR.n136 VGND 0.22037f
C573 VDPWR.n137 VGND 2.55468f
C574 VDPWR.n138 VGND 0.04093f
C575 VDPWR.n139 VGND 0.04093f
C576 VDPWR.n140 VGND 0.10617f
C577 VDPWR.n141 VGND 0.11454f
C578 VDPWR.n142 VGND 0.01488f
C579 VDPWR.n143 VGND 0.21915f
C580 VDPWR.n144 VGND 2.55468f
C581 VDPWR.n145 VGND 0.04899f
C582 VDPWR.n146 VGND 0.04093f
C583 VDPWR.n147 VGND 0.04093f
C584 VDPWR.n148 VGND 0.67366f
C585 VDPWR.n149 VGND 0.01488f
C586 VDPWR.n150 VGND 0.21915f
C587 VDPWR.n151 VGND 0.04879f
C588 VDPWR.n152 VGND 0.04078f
C589 VDPWR.n153 VGND 1.79597f
C590 VDPWR.n154 VGND 0.04092f
C591 VDPWR.n155 VGND 0.04092f
C592 VDPWR.n156 VGND 2.52976f
C593 VDPWR.n157 VGND 0.04879f
C594 VDPWR.n158 VGND 0.04078f
C595 VDPWR.n159 VGND 0.21915f
C596 VDPWR.n160 VGND 0.01488f
C597 VDPWR.n161 VGND 0.22037f
C598 VDPWR.n162 VGND 2.566f
C599 VDPWR.n163 VGND 0.04093f
C600 VDPWR.n164 VGND 0.04168f
C601 VDPWR.n165 VGND 0.04101f
C602 VDPWR.n166 VGND 0.04101f
C603 VDPWR.n167 VGND 0.10639f
C604 VDPWR.n168 VGND 0.04168f
C605 VDPWR.n169 VGND 0.35922f
C606 VDPWR.n170 VGND -0.08114f
C607 VDPWR.n171 VGND 0.03579f
C608 VDPWR.n172 VGND 0.00663f
C609 VDPWR.n173 VGND 0.03176f
C610 VDPWR.n174 VGND 0.10394f
C611 VDPWR.n175 VGND 0.00663f
C612 VDPWR.n176 VGND 0.65798f
C613 VDPWR.n177 VGND 0.20856f
C614 VDPWR.n178 VGND 0.03166f
C615 VDPWR.n179 VGND 0.03176f
C616 VDPWR.n180 VGND 0.02932f
C617 VDPWR.n181 VGND 0.0175f
C618 VDPWR.n182 VGND 0.67992f
C619 VDPWR.n183 VGND 0.39028f
C620 VDPWR.n184 VGND 0.0175f
C621 VDPWR.n185 VGND 0.21034f
C622 VDPWR.n186 VGND 0.03166f
C623 VDPWR.n187 VGND 0.03166f
C624 VDPWR.n188 VGND 0.10394f
C625 VDPWR.n189 VGND 0.67366f
C626 VDPWR.n190 VGND 0.37059f
C627 VDPWR.n191 VGND 0.0058f
C628 VDPWR.n192 VGND 0.10692f
C629 VDPWR.n193 VGND 0.04168f
C630 VDPWR.n194 VGND 0.01921f
C631 VDPWR.n195 VGND 0.03176f
C632 VDPWR.n196 VGND 0.35922f
C633 VDPWR.n197 VGND 0.65798f
C634 VDPWR.n198 VGND 0.02932f
C635 VDPWR.n199 VGND 0.20856f
C636 VDPWR.n200 VGND 2.08134f
C637 VDPWR.n201 VGND 2.45276f
C638 VDPWR.n202 VGND 0.03579f
C639 VDPWR.n203 VGND 0.03176f
C640 VDPWR.n204 VGND 0.11146f
C641 VDPWR.n205 VGND -0.08114f
C642 VDPWR.n206 VGND 0.04101f
C643 VDPWR.n207 VGND 0.04078f
C644 VDPWR.n208 VGND 0.01488f
C645 VDPWR.n209 VGND 0.00663f
C646 VDPWR.n210 VGND 0.00663f
C647 VDPWR.n211 VGND 0.04078f
C648 VDPWR.n212 VGND 0.01488f
C649 VDPWR.n213 VGND 2.23761f
C650 VDPWR.n214 VGND 2.18778f
C651 VDPWR.n215 VGND 0.04101f
C652 VDPWR.n216 VGND 0.10617f
C653 VDPWR.n217 VGND 0.11454f
C654 VDPWR.n218 VGND 0.11558f
C655 VDPWR.n219 VGND 0.10639f
C656 VDPWR.n220 VGND 0.03176f
C657 VDPWR.n221 VGND 0.03579f
C658 VDPWR.n222 VGND 0.03176f
C659 VDPWR.n223 VGND 0.02928f
C660 VDPWR.n224 VGND 0.01417f
C661 VDPWR.n225 VGND 0.02335f
C662 VDPWR.n226 VGND 0.01417f
C663 VDPWR.n227 VGND 0.02928f
C664 VDPWR.n228 VGND 0.21034f
C665 VDPWR.n229 VGND 0.03579f
C666 VDPWR.n230 VGND 0.03176f
C667 VDPWR.n231 VGND 0.03166f
C668 VDPWR.n232 VGND 0.03176f
C669 VDPWR.n233 VGND 0.11146f
C670 VDPWR.n234 VGND 0.01921f
C671 VDPWR.n235 VGND 0.10692f
C672 VDPWR.n236 VGND 0.10617f
C673 VDPWR.n237 VGND 0.11454f
C674 VDPWR.n238 VGND 0.11558f
C675 VDPWR.n239 VGND 0.0058f
C676 VDPWR.n240 VGND 0.37059f
C677 VDPWR.n241 VGND 0.04168f
C678 VDPWR.n242 VGND 1.80956f
C679 VDPWR.n243 VGND 0.40313f
C680 VDPWR.n244 VGND 0.04093f
C681 VDPWR.n245 VGND 0.03761f
C682 VDPWR.n246 VGND 0.04078f
C683 VDPWR.n247 VGND 0.03762f
C684 VDPWR.n248 VGND 0.04092f
C685 VDPWR.n249 VGND 0.50278f
C686 VDPWR.n250 VGND 0.04092f
C687 VDPWR.n251 VGND 0.03762f
C688 VDPWR.n252 VGND 0.04078f
C689 VDPWR.n253 VGND 0.03761f
C690 VDPWR.n254 VGND 0.22037f
C691 VDPWR.n255 VGND 0.04899f
C692 VDPWR.n256 VGND 2.67471f
C693 VDPWR.n257 VGND 0.04092f
C694 VDPWR.n258 VGND 0.04092f
C695 VDPWR.n259 VGND 0.03761f
C696 VDPWR.n260 VGND 0.04078f
C697 VDPWR.n261 VGND 0.01488f
C698 VDPWR.n262 VGND 0.01488f
C699 VDPWR.n263 VGND 0.04078f
C700 VDPWR.n264 VGND 0.03762f
C701 VDPWR.n265 VGND 0.21915f
C702 VDPWR.n266 VGND 0.04879f
C703 VDPWR.n267 VGND 2.67245f
C704 VDPWR.n268 VGND 0.04879f
C705 VDPWR.n269 VGND 0.04092f
C706 VDPWR.n270 VGND 0.04078f
C707 VDPWR.n271 VGND 0.01488f
C708 VDPWR.n272 VGND 0.04078f
C709 VDPWR.n273 VGND 0.04092f
C710 VDPWR.n274 VGND 0.03762f
C711 VDPWR.n275 VGND 0.04078f
C712 VDPWR.n276 VGND 0.03761f
C713 VDPWR.n277 VGND 0.02928f
C714 VDPWR.n278 VGND 0.21034f
C715 VDPWR.n279 VGND 0.0058f
C716 VDPWR.n280 VGND 0.04168f
C717 VDPWR.n281 VGND 1.80956f
C718 VDPWR.n282 VGND 0.04168f
C719 VDPWR.n283 VGND 0.37059f
C720 VDPWR.n284 VGND 0.67366f
C721 VDPWR.n285 VGND 0.22037f
C722 VDPWR.n286 VGND 0.04899f
C723 VDPWR.n287 VGND 2.07907f
C724 VDPWR.n288 VGND 0.04899f
C725 VDPWR.n289 VGND 0.04093f
C726 VDPWR.n290 VGND 0.0058f
C727 VDPWR.n291 VGND 0.11558f
C728 VDPWR.n292 VGND 0.10639f
C729 VDPWR.n293 VGND 0.03166f
C730 VDPWR.n294 VGND 0.00663f
C731 VDPWR.n295 VGND 0.00663f
C732 VDPWR.n296 VGND 0.10394f
C733 VDPWR.n297 VGND -0.08114f
C734 VDPWR.n298 VGND 0.11146f
C735 VDPWR.n299 VGND 0.01921f
C736 VDPWR.n300 VGND 0.35922f
C737 VDPWR.n301 VGND 0.04168f
C738 VDPWR.n302 VGND 1.79597f
C739 VDPWR.n303 VGND 0.04168f
C740 VDPWR.n304 VGND 0.35922f
C741 VDPWR.n305 VGND 0.01921f
C742 VDPWR.n306 VGND 0.11146f
C743 VDPWR.n307 VGND 0.03176f
C744 VDPWR.n308 VGND 2.52976f
C745 VDPWR.n309 VGND 0.03176f
C746 VDPWR.n310 VGND 0.03166f
C747 VDPWR.n311 VGND 0.00663f
C748 VDPWR.n312 VGND 0.00663f
C749 VDPWR.n313 VGND 0.10394f
C750 VDPWR.n314 VGND 0.10639f
C751 VDPWR.n315 VGND 0.03176f
C752 VDPWR.n316 VGND 2.566f
C753 VDPWR.n317 VGND 0.03176f
C754 VDPWR.n318 VGND 0.02928f
C755 VDPWR.n319 VGND 0.01417f
C756 VDPWR.n320 VGND 0.02335f
C757 VDPWR.n321 VGND 0.67992f
C758 VDPWR.n322 VGND 0.5157f
C759 VDPWR.n323 VGND 3.01633f
C760 VDPWR.n324 VGND 0.18492f
C761 VDPWR.n325 VGND 0.14034f
C762 VDPWR.n326 VGND 0.12147f
C763 VDPWR.n327 VGND 0.21068f
C764 VDPWR.n328 VGND 0.40385f
C765 VDPWR.n329 VGND 0.55981f
C766 VDPWR.n330 VGND 0.0175f
C767 VDPWR.n331 VGND 0.21034f
C768 VDPWR.n332 VGND 0.03166f
C769 VDPWR.n333 VGND 0.03579f
C770 VDPWR.n334 VGND 1.1188f
C771 VDPWR.n335 VGND 0.03176f
C772 VDPWR.n336 VGND 0.04093f
C773 VDPWR.n337 VGND 0.90478f
C774 VDPWR.n338 VGND 0.04078f
C775 VDPWR.n339 VGND 1.38506f
C776 VDPWR.n340 VGND 0.9808f
C777 VDPWR.n341 VGND 0.11558f
C778 VDPWR.n342 VGND 0.67366f
C779 VDPWR.n343 VGND 0.04101f
C780 VDPWR.n344 VGND 0.04168f
C781 VDPWR.n345 VGND 0.10617f
C782 VDPWR.n346 VGND 0.25139f
C783 VDPWR.n347 VGND 0.03176f
C784 VDPWR.n348 VGND 0.03579f
C785 VDPWR.n349 VGND 0.21915f
C786 VDPWR.n350 VGND 0.04078f
C787 VDPWR.n351 VGND 0.22037f
C788 VDPWR.n352 VGND 0.03761f
C789 VDPWR.n353 VGND 0.11454f
C790 VDPWR.n354 VGND 0.01488f
C791 VDPWR.n355 VGND 0.01488f
C792 VDPWR.n356 VGND 0.04078f
C793 VDPWR.n357 VGND 0.03762f
C794 VDPWR.n358 VGND 0.04092f
C795 VDPWR.n359 VGND 1.27734f
C796 VDPWR.n360 VGND 0.04093f
C797 VDPWR.n361 VGND 0.04093f
C798 VDPWR.n362 VGND 0.67366f
C799 VDPWR.n363 VGND 0.01488f
C800 VDPWR.n364 VGND 0.21915f
C801 VDPWR.n365 VGND 0.98133f
C802 VDPWR.n366 VGND 0.04078f
C803 VDPWR.n367 VGND 0.89799f
C804 VDPWR.n368 VGND 0.04092f
C805 VDPWR.n369 VGND 0.03176f
C806 VDPWR.n370 VGND 1.09389f
C807 VDPWR.n371 VGND 1.33451f
C808 VDPWR.n372 VGND 0.03579f
C809 VDPWR.n373 VGND 0.03166f
C810 VDPWR.n374 VGND 0.20856f
C811 VDPWR.n375 VGND 0.00663f
C812 VDPWR.n376 VGND 0.21034f
C813 VDPWR.n377 VGND 0.03579f
C814 VDPWR.n378 VGND 0.04078f
C815 VDPWR.n379 VGND 0.01488f
C816 VDPWR.n380 VGND 1.1188f
C817 VDPWR.n381 VGND 0.00663f
C818 VDPWR.n382 VGND 0.03166f
C819 VDPWR.n383 VGND 0.03176f
C820 VDPWR.n384 VGND 0.04101f
C821 VDPWR.n385 VGND 0.04101f
C822 VDPWR.n386 VGND 0.10639f
C823 VDPWR.n387 VGND 0.65798f
C824 VDPWR.n388 VGND 0.04168f
C825 VDPWR.n389 VGND 0.35922f
C826 VDPWR.n390 VGND 0.10394f
C827 VDPWR.n391 VGND -0.08114f
C828 VDPWR.n392 VGND 0.11146f
C829 VDPWR.n393 VGND 0.01921f
C830 VDPWR.n394 VGND 0.10692f
C831 VDPWR.n395 VGND 0.10617f
C832 VDPWR.n396 VGND 0.11454f
C833 VDPWR.n397 VGND 0.11558f
C834 VDPWR.n398 VGND 0.0058f
C835 VDPWR.n399 VGND 0.37059f
C836 VDPWR.n400 VGND 0.04168f
C837 VDPWR.n401 VGND 0.90478f
C838 VDPWR.n402 VGND 0.20157f
C839 VDPWR.n403 VGND 1.283f
C840 VDPWR.n404 VGND 0.03176f
C841 VDPWR.n405 VGND 0.02928f
C842 VDPWR.n406 VGND 0.73645f
C843 VDPWR.n407 VGND 0.79274f
C844 VDPWR.n408 VGND 1.76097f
C845 VDPWR.n409 VGND 0.28953f
C846 VDPWR.n410 VGND 0.40361f
C847 VDPWR.n411 VGND 0.55981f
C848 VDPWR.n412 VGND 0.04332f
C849 VDPWR.n413 VGND 0.01417f
C850 VDPWR.n414 VGND 0.0175f
C851 VDPWR.n415 VGND 0.02932f
C852 VDPWR.n416 VGND 0.03176f
C853 VDPWR.n417 VGND 1.26488f
C854 VDPWR.n418 VGND 0.25139f
C855 VDPWR.n419 VGND 0.04092f
C856 VDPWR.n420 VGND 0.03762f
C857 VDPWR.n421 VGND 0.04078f
C858 VDPWR.n422 VGND 0.03761f
C859 VDPWR.n423 VGND 0.22037f
C860 VDPWR.n424 VGND 0.04899f
C861 VDPWR.n425 VGND 1.33736f
C862 VDPWR.n426 VGND 0.89799f
C863 VDPWR.n427 VGND 1.22638f
C864 VDPWR.n428 VGND 1.33622f
C865 VDPWR.n429 VGND 0.04879f
C866 VDPWR.n430 VGND 0.04092f
C867 VDPWR.n431 VGND 0.10692f
C868 VDPWR.n432 VGND 0.10639f
C869 VDPWR.n433 VGND 0.03166f
C870 VDPWR.n434 VGND 0.00663f
C871 VDPWR.n435 VGND 0.00663f
C872 VDPWR.n436 VGND 0.10394f
C873 VDPWR.n437 VGND -0.08114f
C874 VDPWR.n438 VGND 0.11146f
C875 VDPWR.n439 VGND 0.01921f
C876 VDPWR.n440 VGND 0.35922f
C877 VDPWR.n441 VGND 0.65798f
C878 VDPWR.n442 VGND 0.20856f
C879 VDPWR.n443 VGND 0.02932f
C880 VDPWR.n444 VGND 0.03176f
C881 VDPWR.n445 VGND 1.26488f
C882 VDPWR.n446 VGND 1.09389f
C883 VDPWR.n447 VGND 0.04101f
C884 VDPWR.n448 VGND 0.04168f
C885 VDPWR.n449 VGND 0.37059f
C886 VDPWR.n450 VGND 0.0058f
C887 VDPWR.n451 VGND 0.04093f
C888 VDPWR.n452 VGND 0.20157f
C889 VDPWR.n453 VGND 1.283f
C890 VDPWR.n454 VGND 0.03176f
C891 VDPWR.n455 VGND 0.02928f
C892 VDPWR.n456 VGND 0.01417f
C893 VDPWR.n457 VGND 0.04332f
C894 VDPWR.n458 VGND 0.73645f
C895 VDPWR.n459 VGND 0.79274f
C896 VDPWR.n460 VGND 2.00086f
C897 VDPWR.n461 VGND 0.15589f
C898 VDPWR.n462 VGND 1.14196f
C899 VDPWR.n463 VGND 1.99709f
C900 VDPWR.n464 VGND 1.15985f
C901 VDPWR.n465 VGND 2.69328f
C902 VDPWR.n466 VGND 3.53752f
C903 VDPWR.n467 VGND 3.627f
C904 VDPWR.n468 VGND 3.90883f
C905 VDPWR.n469 VGND 0.00544f
C906 VDPWR.n470 VGND 0.10808f
C907 VDPWR.n471 VGND 0.0078f
C908 VDPWR.n472 VGND 0.01556f
C909 VDPWR.n473 VGND 0.01556f
C910 VDPWR.n474 VGND 0.7724f
C911 VDPWR.n475 VGND 0.01519f
C912 VDPWR.n476 VGND 0.7724f
C913 VDPWR.n477 VGND 0.01519f
C914 VDPWR.n478 VGND 0.01519f
C915 VDPWR.n479 VGND 0.01556f
C916 VDPWR.n480 VGND 0.01556f
C917 VDPWR.n481 VGND 0.01517f
C918 VDPWR.n482 VGND 0.0078f
C919 VDPWR.n483 VGND 0.01556f
C920 VDPWR.n484 VGND 0.01556f
C921 VDPWR.n485 VGND 0.7724f
C922 VDPWR.n486 VGND 0.01519f
C923 VDPWR.n487 VGND 0.01519f
C924 VDPWR.n488 VGND 0.01519f
C925 VDPWR.n489 VGND 0.7724f
C926 VDPWR.n490 VGND 0.01556f
C927 VDPWR.n491 VGND 0.01556f
C928 VDPWR.n492 VGND 0.0078f
C929 VDPWR.n493 VGND 0.01519f
C930 VDPWR.n494 VGND 0.01517f
C931 VDPWR.n495 VGND 0.01519f
C932 VDPWR.n496 VGND 1.19788f
C933 VDPWR.n497 VGND 0.01519f
C934 VDPWR.n498 VGND 0.01517f
C935 VDPWR.n499 VGND 0.00544f
C936 VDPWR.n500 VGND 0.10808f
C937 VDPWR.n501 VGND 0.02417f
C938 VDPWR.n502 VGND 0.00544f
C939 VDPWR.n503 VGND 0.0078f
C940 VDPWR.n504 VGND 0.01519f
C941 VDPWR.n505 VGND 0.01519f
C942 VDPWR.n506 VGND 1.19788f
C943 VDPWR.n507 VGND 0.01519f
C944 VDPWR.n508 VGND 0.01517f
C945 VDPWR.n509 VGND 0.00544f
C946 VDPWR.n510 VGND 0.12217f
C947 VDPWR.n511 VGND 0.66392f
C948 VDPWR.n512 VGND 1.18771f
C949 VDPWR.n513 VGND 0.65572f
C950 VDPWR.n514 VGND 3.65583f
C951 VDPWR.n515 VGND 1.74868f
C952 VDPWR.n516 VGND 0.77946f
C953 VDPWR.n517 VGND 0.00544f
C954 VDPWR.n518 VGND 0.10808f
C955 VDPWR.n519 VGND 0.0078f
C956 VDPWR.n520 VGND 0.01556f
C957 VDPWR.n521 VGND 0.01556f
C958 VDPWR.n522 VGND 0.7724f
C959 VDPWR.n523 VGND 0.01519f
C960 VDPWR.n524 VGND 0.7724f
C961 VDPWR.n525 VGND 0.01519f
C962 VDPWR.n526 VGND 0.01519f
C963 VDPWR.n527 VGND 0.01556f
C964 VDPWR.n528 VGND 0.01556f
C965 VDPWR.n529 VGND 0.01517f
C966 VDPWR.n530 VGND 0.0078f
C967 VDPWR.n531 VGND 0.01556f
C968 VDPWR.n532 VGND 0.01556f
C969 VDPWR.n533 VGND 0.7724f
C970 VDPWR.n534 VGND 0.01519f
C971 VDPWR.n535 VGND 0.01519f
C972 VDPWR.n536 VGND 0.01519f
C973 VDPWR.n537 VGND 0.7724f
C974 VDPWR.n538 VGND 0.01556f
C975 VDPWR.n539 VGND 0.01556f
C976 VDPWR.n540 VGND 0.0078f
C977 VDPWR.n541 VGND 0.01519f
C978 VDPWR.n542 VGND 0.01517f
C979 VDPWR.n543 VGND 0.01519f
C980 VDPWR.n544 VGND 1.19788f
C981 VDPWR.n545 VGND 0.01519f
C982 VDPWR.n546 VGND 0.01517f
C983 VDPWR.n547 VGND 0.00544f
C984 VDPWR.n548 VGND 0.10808f
C985 VDPWR.n549 VGND 0.02417f
C986 VDPWR.n550 VGND 0.00544f
C987 VDPWR.n551 VGND 0.0078f
C988 VDPWR.n552 VGND 0.01519f
C989 VDPWR.n553 VGND 0.01519f
C990 VDPWR.n554 VGND 1.19788f
C991 VDPWR.n555 VGND 0.01519f
C992 VDPWR.n556 VGND 0.01517f
C993 VDPWR.n557 VGND 0.00544f
C994 VDPWR.n558 VGND 0.12217f
C995 VDPWR.n559 VGND 0.6651f
C996 VDPWR.n560 VGND 0.71585f
C997 VDPWR.n561 VGND 1.83185f
C998 VDPWR.n562 VGND 3.11219f
C999 VDPWR.n563 VGND 0.59006f
C1000 VDPWR.n564 VGND 0.46406f
C1001 VDPWR.n565 VGND 0.58632f
C1002 VDPWR.n566 VGND 0.0175f
C1003 VDPWR.n567 VGND 0.21034f
C1004 VDPWR.n568 VGND 0.03166f
C1005 VDPWR.n569 VGND 0.03579f
C1006 VDPWR.n570 VGND 1.1188f
C1007 VDPWR.n571 VGND 0.20157f
C1008 VDPWR.n572 VGND 0.03166f
C1009 VDPWR.n573 VGND 0.00663f
C1010 VDPWR.n574 VGND 0.00663f
C1011 VDPWR.n575 VGND 0.10394f
C1012 VDPWR.n576 VGND 0.0058f
C1013 VDPWR.n577 VGND 0.10617f
C1014 VDPWR.n578 VGND 0.04078f
C1015 VDPWR.n579 VGND 0.04078f
C1016 VDPWR.n580 VGND 0.04092f
C1017 VDPWR.n581 VGND 0.04093f
C1018 VDPWR.n582 VGND 0.03761f
C1019 VDPWR.n583 VGND 0.22037f
C1020 VDPWR.n584 VGND 0.04101f
C1021 VDPWR.n585 VGND 0.04168f
C1022 VDPWR.n586 VGND -0.08114f
C1023 VDPWR.n587 VGND 0.25139f
C1024 VDPWR.n588 VGND 0.03176f
C1025 VDPWR.n589 VGND 0.03579f
C1026 VDPWR.n590 VGND 0.10692f
C1027 VDPWR.n591 VGND 0.03762f
C1028 VDPWR.n592 VGND 0.04092f
C1029 VDPWR.n593 VGND 0.89799f
C1030 VDPWR.n594 VGND 1.33451f
C1031 VDPWR.n595 VGND 0.98133f
C1032 VDPWR.n596 VGND 0.21915f
C1033 VDPWR.n597 VGND 0.02932f
C1034 VDPWR.n598 VGND 0.20856f
C1035 VDPWR.n599 VGND 0.65798f
C1036 VDPWR.n600 VGND 0.35922f
C1037 VDPWR.n601 VGND 0.01921f
C1038 VDPWR.n602 VGND 0.11146f
C1039 VDPWR.n603 VGND 0.03176f
C1040 VDPWR.n604 VGND 1.26488f
C1041 VDPWR.n605 VGND 1.09389f
C1042 VDPWR.n606 VGND 0.04101f
C1043 VDPWR.n607 VGND 0.67366f
C1044 VDPWR.n608 VGND 0.37059f
C1045 VDPWR.n609 VGND 0.04168f
C1046 VDPWR.n610 VGND 0.90478f
C1047 VDPWR.n611 VGND 1.27734f
C1048 VDPWR.n612 VGND 0.73703f
C1049 VDPWR.n613 VGND 0.04101f
C1050 VDPWR.n614 VGND 0.04101f
C1051 VDPWR.n615 VGND 0.03738f
C1052 VDPWR.n616 VGND 0.02091f
C1053 VDPWR.n618 VGND 0.47371f
C1054 VDPWR.n619 VGND 0.0229f
C1055 VDPWR.n620 VGND 0.01909f
C1056 VDPWR.n621 VGND 0.65247f
C1057 VDPWR.n622 VGND 0.29316f
C1058 VDPWR.n623 VGND 0.1943f
C1059 VDPWR.n624 VGND 0.1916f
C1060 VDPWR.n625 VGND 0.02322f
C1061 VDPWR.n626 VGND 0.04281f
C1062 VDPWR.n627 VGND 0.04168f
C1063 VDPWR.n628 VGND 1.16281f
C1064 VDPWR.n629 VGND 1.7504f
C1065 VDPWR.n630 VGND 0.04899f
C1066 VDPWR.n631 VGND 0.04093f
C1067 VDPWR.n632 VGND 0.04078f
C1068 VDPWR.n633 VGND 0.01488f
C1069 VDPWR.n634 VGND 0.01488f
C1070 VDPWR.n635 VGND 0.11454f
C1071 VDPWR.n636 VGND 0.11558f
C1072 VDPWR.n637 VGND 0.10639f
C1073 VDPWR.n638 VGND 0.03176f
C1074 VDPWR.n639 VGND 1.283f
C1075 VDPWR.n640 VGND 0.03176f
C1076 VDPWR.n641 VGND 0.02928f
C1077 VDPWR.n642 VGND 0.01417f
C1078 VDPWR.n643 VGND 0.03134f
C1079 VDPWR.n644 VGND 0.42173f
C1080 VDPWR.n645 VGND 0.31943f
C1081 VDPWR.n646 VGND 0.27276f
C1082 VDPWR.n647 VGND 1.61763f
C1083 VDPWR.n648 VGND 1.15456f
C1084 VDPWR.n649 VGND 4.11699f
C1085 VDPWR.n650 VGND 3.51846f
C1086 VDPWR.n651 VGND 10.2621f
C1087 VDPWR.n652 VGND 11.9507f
C1088 VDPWR.n653 VGND 11.3581f
C1089 VDPWR.n654 VGND 10.2806f
C1090 VDPWR.n655 VGND 1.06341f
C1091 VDPWR.n656 VGND 0.44306f
C1092 VDPWR.n657 VGND 0.17671f
C1093 VDPWR.n658 VGND 0.43971f
C1094 VDPWR.n659 VGND 3.24805f
C1095 VDPWR.n660 VGND 2.27041f
C1096 VDPWR.n661 VGND 4.68567f
C1097 VDPWR.n662 VGND 3.12958f
C1098 VDPWR.n663 VGND 3.15083f
C1099 VDPWR.n664 VGND 1.99155f
C1100 VDPWR.n665 VGND 0.00232f
C1101 VDPWR.n666 VGND 0.13616f
C1102 VDPWR.n667 VGND 0.00233f
C1103 VDPWR.n668 VGND 0.01024f
C1104 VDPWR.n669 VGND 0.01519f
C1105 VDPWR.n670 VGND 0.00976f
C1106 VDPWR.n671 VGND 0.01519f
C1107 VDPWR.n672 VGND 0.22856f
C1108 VDPWR.n673 VGND 0.0101f
C1109 VDPWR.n674 VGND 0.01519f
C1110 VDPWR.n675 VGND 0.22856f
C1111 VDPWR.n676 VGND 0.01556f
C1112 VDPWR.n677 VGND 0.01556f
C1113 VDPWR.n678 VGND 0.01517f
C1114 VDPWR.n679 VGND 0.00544f
C1115 VDPWR.n680 VGND 0.00544f
C1116 VDPWR.n681 VGND 0.10808f
C1117 VDPWR.n682 VGND 0.0078f
C1118 VDPWR.n683 VGND 0.01556f
C1119 VDPWR.n684 VGND 0.01556f
C1120 VDPWR.n685 VGND 0.22856f
C1121 VDPWR.n686 VGND 0.01556f
C1122 VDPWR.n687 VGND 0.01556f
C1123 VDPWR.n688 VGND 0.0078f
C1124 VDPWR.n689 VGND 0.01556f
C1125 VDPWR.n690 VGND 0.01556f
C1126 VDPWR.n691 VGND 0.0078f
C1127 VDPWR.n692 VGND 0.01519f
C1128 VDPWR.n693 VGND 0.01517f
C1129 VDPWR.n694 VGND 0.01519f
C1130 VDPWR.n695 VGND 0.01519f
C1131 VDPWR.n696 VGND 0.1895f
C1132 VDPWR.n697 VGND 0.01519f
C1133 VDPWR.n698 VGND 0.01519f
C1134 VDPWR.n699 VGND 0.1895f
C1135 VDPWR.n700 VGND 0.01519f
C1136 VDPWR.n701 VGND 0.01519f
C1137 VDPWR.n702 VGND 0.01517f
C1138 VDPWR.n703 VGND 0.01519f
C1139 VDPWR.n704 VGND 0.19095f
C1140 VDPWR.n705 VGND 0.01519f
C1141 VDPWR.n706 VGND 0.01517f
C1142 VDPWR.n707 VGND 0.00544f
C1143 VDPWR.n708 VGND 0.02417f
C1144 VDPWR.n709 VGND 0.10808f
C1145 VDPWR.n710 VGND 0.0243f
C1146 VDPWR.n711 VGND 0.00544f
C1147 VDPWR.n712 VGND 0.0078f
C1148 VDPWR.n713 VGND 0.01519f
C1149 VDPWR.n714 VGND 0.01519f
C1150 VDPWR.n715 VGND 0.19095f
C1151 VDPWR.n716 VGND 0.19095f
C1152 VDPWR.n717 VGND 0.0101f
C1153 VDPWR.n718 VGND 0.01024f
C1154 VDPWR.n719 VGND 0.00976f
C1155 VDPWR.n720 VGND 0.00976f
C1156 VDPWR.n721 VGND 0.00976f
C1157 VDPWR.n722 VGND 0.22856f
C1158 VDPWR.n723 VGND 0.00464f
C1159 VDPWR.n724 VGND 0.00464f
C1160 VDPWR.n725 VGND 0.00976f
C1161 VDPWR.n726 VGND 0.00976f
C1162 VDPWR.n727 VGND 0.0101f
C1163 VDPWR.n728 VGND 0.00976f
C1164 VDPWR.n729 VGND 0.01024f
C1165 VDPWR.n730 VGND 0.01024f
C1166 VDPWR.n731 VGND 0.00974f
C1167 VDPWR.n732 VGND 0.0101f
C1168 VDPWR.n733 VGND 0.01519f
C1169 VDPWR.n734 VGND 0.01519f
C1170 VDPWR.n735 VGND 0.00976f
C1171 VDPWR.n736 VGND 0.00976f
C1172 VDPWR.n737 VGND 0.01519f
C1173 VDPWR.n738 VGND 0.01519f
C1174 VDPWR.n739 VGND 0.22856f
C1175 VDPWR.n740 VGND 0.0101f
C1176 VDPWR.n741 VGND 0.0101f
C1177 VDPWR.n742 VGND 0.01024f
C1178 VDPWR.n743 VGND 0.00233f
C1179 VDPWR.n744 VGND 0.00544f
C1180 VDPWR.n745 VGND 0.0078f
C1181 VDPWR.n746 VGND 0.01556f
C1182 VDPWR.n747 VGND 0.01556f
C1183 VDPWR.n748 VGND 0.22856f
C1184 VDPWR.n749 VGND 0.01556f
C1185 VDPWR.n750 VGND 0.01556f
C1186 VDPWR.n751 VGND 0.0078f
C1187 VDPWR.n752 VGND 0.22856f
C1188 VDPWR.n753 VGND 0.01519f
C1189 VDPWR.n754 VGND 0.01556f
C1190 VDPWR.n755 VGND 0.01556f
C1191 VDPWR.n756 VGND 0.00544f
C1192 VDPWR.n757 VGND 0.0078f
C1193 VDPWR.n758 VGND 0.01556f
C1194 VDPWR.n759 VGND 0.01556f
C1195 VDPWR.n760 VGND 0.01517f
C1196 VDPWR.n761 VGND 0.10808f
C1197 VDPWR.n762 VGND 0.03894f
C1198 VDPWR.n763 VGND 0.00544f
C1199 VDPWR.n764 VGND 0.0078f
C1200 VDPWR.n765 VGND 0.01519f
C1201 VDPWR.n766 VGND 0.01519f
C1202 VDPWR.n767 VGND 0.19095f
C1203 VDPWR.n768 VGND 0.01519f
C1204 VDPWR.n769 VGND 0.01519f
C1205 VDPWR.n770 VGND 0.01517f
C1206 VDPWR.n771 VGND 0.01519f
C1207 VDPWR.n772 VGND 0.1895f
C1208 VDPWR.n773 VGND 0.01519f
C1209 VDPWR.n774 VGND 0.01519f
C1210 VDPWR.n775 VGND 0.1895f
C1211 VDPWR.n776 VGND 0.01519f
C1212 VDPWR.n777 VGND 0.01519f
C1213 VDPWR.n778 VGND 0.01517f
C1214 VDPWR.n779 VGND 0.01519f
C1215 VDPWR.n780 VGND 0.22856f
C1216 VDPWR.n781 VGND 0.0101f
C1217 VDPWR.n782 VGND 0.0101f
C1218 VDPWR.n783 VGND 0.00976f
C1219 VDPWR.n784 VGND 0.00976f
C1220 VDPWR.n785 VGND 0.00976f
C1221 VDPWR.n786 VGND 0.00464f
C1222 VDPWR.n787 VGND 0.22856f
C1223 VDPWR.n788 VGND 0.00976f
C1224 VDPWR.n789 VGND 0.01024f
C1225 VDPWR.n790 VGND 0.00976f
C1226 VDPWR.n791 VGND 0.00976f
C1227 VDPWR.n792 VGND 0.00464f
C1228 VDPWR.n793 VGND 0.22856f
C1229 VDPWR.n794 VGND 0.22856f
C1230 VDPWR.n795 VGND 0.01024f
C1231 VDPWR.n796 VGND 0.01024f
C1232 VDPWR.n797 VGND 0.00976f
C1233 VDPWR.n798 VGND 0.0101f
C1234 VDPWR.n799 VGND 0.01519f
C1235 VDPWR.n800 VGND 0.01519f
C1236 VDPWR.n801 VGND 0.19095f
C1237 VDPWR.n802 VGND 0.19095f
C1238 VDPWR.n803 VGND 0.01519f
C1239 VDPWR.n804 VGND 0.01517f
C1240 VDPWR.n805 VGND 0.00544f
C1241 VDPWR.n806 VGND 0.02417f
C1242 VDPWR.n807 VGND 0.10808f
C1243 VDPWR.n808 VGND 0.08624f
C1244 VDPWR.n809 VGND 0.06829f
C1245 VDPWR.n810 VGND 0.00232f
C1246 VDPWR.n811 VGND 0.00974f
C1247 VDPWR.n812 VGND 0.0101f
C1248 VDPWR.n813 VGND 0.01519f
C1249 VDPWR.n814 VGND 0.01519f
C1250 VDPWR.n815 VGND 0.19095f
C1251 VDPWR.n816 VGND 0.19095f
C1252 VDPWR.n817 VGND 0.0101f
C1253 VDPWR.n818 VGND 0.0101f
C1254 VDPWR.n819 VGND 0.01519f
C1255 VDPWR.n820 VGND 0.00976f
C1256 VDPWR.n821 VGND 0.01024f
C1257 VDPWR.n822 VGND 0.01024f
C1258 VDPWR.n823 VGND 0.00976f
C1259 VDPWR.n824 VGND 0.0101f
C1260 VDPWR.n825 VGND 0.01519f
C1261 VDPWR.n826 VGND 0.0101f
C1262 VDPWR.n827 VGND 0.22856f
C1263 VDPWR.n828 VGND 0.0101f
C1264 VDPWR.n829 VGND 0.00976f
C1265 VDPWR.n830 VGND 0.01024f
C1266 VDPWR.n831 VGND 0.01024f
C1267 VDPWR.n832 VGND 0.00976f
C1268 VDPWR.n833 VGND 0.00233f
C1269 VDPWR.n834 VGND 0.00464f
C1270 VDPWR.n835 VGND 0.22856f
C1271 VDPWR.n836 VGND 0.00464f
C1272 VDPWR.n837 VGND 0.00976f
C1273 VDPWR.n838 VGND 0.0101f
C1274 VDPWR.n839 VGND 0.22856f
C1275 VDPWR.n840 VGND 0.0101f
C1276 VDPWR.n841 VGND 0.0101f
C1277 VDPWR.n842 VGND 0.00974f
C1278 VDPWR.n843 VGND 0.00232f
C1279 VDPWR.n844 VGND 0.06808f
C1280 VDPWR.n845 VGND 0.03646f
C1281 VDPWR.n846 VGND 0.36028f
C1282 VDPWR.n847 VGND 0.29699f
C1283 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A VGND 0.74657f
C1284 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G VGND 0.61957f
C1285 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin VGND 0.52606f
C1286 uo_out[2] VGND 3.31864f
C1287 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin VGND 0.52606f
C1288 uo_out[1] VGND 1.91344f
C1289 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin VGND 0.52752f
C1290 uo_out[0] VGND 1.64603f
C1291 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin VGND 0.52606f
C1292 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out VGND 1.20912f
C1293 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin VGND 0.52707f
C1294 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out VGND 1.2937f
C1295 VDPWR VGND 0.45752p
C1296 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin VGND 0.54717f
C1297 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out VGND 1.40293f
C1298 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin VGND 0.52756f
C1299 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 VGND 0.22292f
C1300 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin VGND 0.52606f
C1301 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out VGND 0.28552f
C1302 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin VGND 0.52645f
C1303 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out VGND 0.30478f
C1304 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin VGND 0.53627f
C1305 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out VGND 0.45287f
C1306 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/m1_n100_n100# VGND 0.10852f
C1307 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VGND 1.29945f
C1308 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in VGND 0.81081f
C1309 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G VGND 0.55523f
C1310 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VGND 3.05907f
C1311 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B VGND 0.42095f
C1312 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G VGND 0.55051f
C1313 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G VGND 0.5548f
C1314 ua[0] VGND 69.92041f
C1315 flashADC_3bit_0/comp_p_6/tail VGND 1.94675f
C1316 uio_out[1] VGND 12.2039f
C1317 flashADC_3bit_0/comp_p_6/latch_right VGND 3.82409f
C1318 flashADC_3bit_0/comp_p_6/out_left VGND 2.23346f
C1319 flashADC_3bit_0/comp_p_6/latch_left VGND 10.96687f
C1320 flashADC_3bit_0/comp_p_5/tail VGND 1.09616f
C1321 uio_out[0] VGND 14.97629f
C1322 flashADC_3bit_0/comp_p_5/latch_right VGND 3.4916f
C1323 flashADC_3bit_0/comp_p_5/out_left VGND 3.34218f
C1324 flashADC_3bit_0/comp_p_5/latch_left VGND 3.68553f
C1325 flashADC_3bit_0/comp_p_4/tail VGND 1.09616f
C1326 uo_out[7] VGND 12.03439f
C1327 flashADC_3bit_0/comp_p_4/latch_right VGND 3.4916f
C1328 flashADC_3bit_0/comp_p_4/out_left VGND 2.12858f
C1329 flashADC_3bit_0/comp_p_4/latch_left VGND 9.16368f
C1330 flashADC_3bit_0/comp_p_3/tail VGND 1.46483f
C1331 uo_out[6] VGND 10.30018f
C1332 flashADC_3bit_0/comp_p_3/latch_right VGND 3.54536f
C1333 flashADC_3bit_0/comp_p_3/out_left VGND 2.61512f
C1334 flashADC_3bit_0/comp_p_3/latch_left VGND 3.73577f
C1335 flashADC_3bit_0/comp_p_2/tail VGND 1.42426f
C1336 uo_out[5] VGND 9.89908f
C1337 flashADC_3bit_0/comp_p_2/latch_right VGND 3.52097f
C1338 flashADC_3bit_0/comp_p_2/out_left VGND 2.45831f
C1339 flashADC_3bit_0/comp_p_2/latch_left VGND 9.18686f
C1340 flashADC_3bit_0/comp_p_0/tail VGND 1.18403f
C1341 uo_out[4] VGND 8.01901f
C1342 flashADC_3bit_0/comp_p_0/latch_right VGND 10.84439f
C1343 flashADC_3bit_0/comp_p_0/out_left VGND 3.21577f
C1344 flashADC_3bit_0/comp_p_0/latch_left VGND 3.69778f
C1345 flashADC_3bit_0/comp_p_1/tail VGND 1.19602f
C1346 uo_out[3] VGND 7.65664f
C1347 flashADC_3bit_0/comp_p_1/latch_right VGND 3.50878f
C1348 flashADC_3bit_0/comp_p_1/out_left VGND 3.65291f
C1349 flashADC_3bit_0/comp_p_1/latch_left VGND 3.70233f
C1350 flashADC_3bit_0/comp_p_0/vinn VGND 5.35191f
C1351 flashADC_3bit_0/comp_p_2/vinn VGND 4.33268f
C1352 flashADC_3bit_0/comp_p_3/vinn VGND 7.55153f
C1353 flashADC_3bit_0/comp_p_4/vinn VGND 3.99482f
C1354 flashADC_3bit_0/comp_p_5/vinn VGND 4.91936f
C1355 flashADC_3bit_0/comp_p_6/vinn VGND 7.43265f
C1356 flashADC_3bit_0/comp_p_1/vinn VGND 6.00724f
C1357 ua[1] VGND 26.34101f
C1358 flashADC_3bit_0/vbias_generation_0/bias_n VGND 2.13825f
C1359 flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 VGND 1.69696f
C1360 flashADC_3bit_0/vbias_generation_0/XR_bias_3/R2 VGND 1.58093f
C1361 flashADC_3bit_0/vbias_generation_0/XR_bias_2/R2 VGND 1.64787f
C1362 flashADC_3bit_0/comp_p_6/vbias_p VGND 13.60684f
.ends

