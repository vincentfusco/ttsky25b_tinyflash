* NGSPICE file created from flashADC_3bit_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9 B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_1p41 l=7
C0 R2 R1 0.01325f
C1 R2 B 0.82332f
C2 R1 B 0.82332f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ELBHUY B D S G
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 D G 0.11229f
C1 S G 0.11229f
C2 S D 0.27388f
C3 S B 0.59197f
C4 D B 0.59197f
C5 G B 0.75059f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_VTBKAA B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 S G 0.21915f
C1 D S 0.54671f
C2 G B 0.43443f
C3 D B 0.634f
C4 S B 0.634f
C5 D G 0.21915f
C6 S VSUBS 0.51455f
C7 D VSUBS 0.51455f
C8 G VSUBS 0.36418f
C9 B VSUBS 5.72384f
.ends

.subckt vbias_generation bias_n vdd XR_bias_2/R2 XR_bias_4/R1 XR_bias_3/R2 bias_p
+ vss
XXR_bias_1 vss XR_bias_2/R2 bias_p sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_2 vss XR_bias_3/R2 XR_bias_2/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_3 vss XR_bias_4/R1 XR_bias_3/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_4 vss XR_bias_4/R1 bias_n sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXMn_bias vss bias_n vss bias_n sky130_fd_pr__nfet_01v8_lvt_ELBHUY
XXMp_bias vdd bias_p vdd bias_p vss sky130_fd_pr__pfet_01v8_lvt_VTBKAA
C0 XR_bias_3/R2 XR_bias_2/R2 0
C1 XR_bias_4/R1 XR_bias_2/R2 0.06887f
C2 bias_p XR_bias_2/R2 0.05112f
C3 bias_n XR_bias_3/R2 0.06908f
C4 bias_n XR_bias_4/R1 0
C5 bias_p vdd 0.22745f
C6 XR_bias_4/R1 XR_bias_3/R2 0
C7 bias_p XR_bias_3/R2 0.06932f
C8 bias_p XR_bias_4/R1 0
C9 XR_bias_2/R2 vdd 0.01866f
C10 vdd vss 6.78775f
C11 bias_n vss 2.48381f
C12 XR_bias_4/R1 vss 1.63605f
C13 XR_bias_3/R2 vss 1.57785f
C14 XR_bias_2/R2 vss 1.57097f
C15 bias_p vss 1.64123f
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_JT48NU B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_5p73 l=5.73
C0 R2 R1 0.06813f
C1 R2 B 1.74197f
C2 R1 B 1.74197f
.ends

.subckt res_ladder_vref ref2 ref5 ref6 vref ref3 ref1 ref0 ref4 vss
XXR1 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR2 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR10 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR3 vss ref6 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR4 vss ref4 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR5 vss ref4 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR6 vss ref2 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR7 vss ref2 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR8 vss ref0 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR9 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
C0 ref5 ref4 0
C1 ref3 ref2 0
C2 ref3 ref5 0.06887f
C3 ref3 ref1 0.06887f
C4 ref0 ref2 0.06887f
C5 ref3 ref4 0
C6 ref6 ref5 0
C7 ref6 vref 0.16095f
C8 ref2 ref1 0
C9 vref ref5 0.06887f
C10 ref2 ref4 0.06887f
C11 ref6 ref4 0.06887f
C12 ref0 ref1 0
C13 ref1 vss 3.4889f
C14 ref2 vss 3.42003f
C15 ref3 vss 3.42003f
C16 ref4 vss 3.42003f
C17 ref5 vss 3.42003f
C18 ref6 vss 5.161f
C19 ref0 vss 5.32418f
C20 vref vss 4.57377f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MMMA4V a_n260_n698# a_100_n500# a_n158_n500# a_n100_n588#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n698# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 a_n100_n588# a_n158_n500# 0.11229f
C1 a_n100_n588# a_100_n500# 0.11229f
C2 a_n158_n500# a_100_n500# 0.27388f
C3 a_100_n500# a_n260_n698# 0.5905f
C4 a_n158_n500# a_n260_n698# 0.5905f
C5 a_n100_n588# a_n260_n698# 0.7183f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_5VNMZ8 a_n100_n897# a_100_n800# w_n296_n1019#
+ a_n158_n800# VSUBS
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n296_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
C0 w_n296_n1019# a_n100_n897# 0.43443f
C1 a_100_n800# a_n158_n800# 0.43758f
C2 w_n296_n1019# a_100_n800# 0.51205f
C3 a_n100_n897# a_100_n800# 0.17641f
C4 w_n296_n1019# a_n158_n800# 0.51205f
C5 a_n100_n897# a_n158_n800# 0.17641f
C6 a_100_n800# VSUBS 0.41369f
C7 a_n158_n800# VSUBS 0.41369f
C8 a_n100_n897# VSUBS 0.36418f
C9 w_n296_n1019# VSUBS 4.82082f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHMAL2 a_n260_n574# a_100_n400# a_n158_n400# a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n260_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
C0 a_n100_n488# a_n158_n400# 0.09092f
C1 a_n100_n488# a_100_n400# 0.09092f
C2 a_n158_n400# a_100_n400# 0.21931f
C3 a_100_n400# a_n260_n574# 0.48057f
C4 a_n158_n400# a_n260_n574# 0.48057f
C5 a_n100_n488# a_n260_n574# 0.74751f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GUWLND a_n158_n1000# a_n100_n1097# w_n296_n1219#
+ a_100_n1000# VSUBS
X0 a_100_n1000# a_n100_n1097# a_n158_n1000# w_n296_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 w_n296_n1219# a_n100_n1097# 0.43443f
C1 a_100_n1000# a_n158_n1000# 0.54671f
C2 w_n296_n1219# a_100_n1000# 0.634f
C3 a_n100_n1097# a_100_n1000# 0.21915f
C4 w_n296_n1219# a_n158_n1000# 0.634f
C5 a_n100_n1097# a_n158_n1000# 0.21915f
C6 a_100_n1000# VSUBS 0.51455f
C7 a_n158_n1000# VSUBS 0.51455f
C8 a_n100_n1097# VSUBS 0.36418f
C9 w_n296_n1219# VSUBS 5.72384f
.ends

.subckt comp_p vinp vinn vbias_p vdd tail vout latch_right out_left latch_left vss
XXMn_cs_left vss latch_right vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_out out_left vdd vdd vout vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_diode_left1 vss latch_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_AHMAL2
XXMn_cs_right1 vss latch_left vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_diode_right vss latch_right vss latch_right sky130_fd_pr__nfet_01v8_lvt_AHMAL2
Xsky130_fd_pr__pfet_01v8_lvt_5VNMZ8_0 out_left vdd vdd out_left vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_out_left vss out_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_out_right vss vout vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_tail tail vbias_p vdd vdd vss sky130_fd_pr__pfet_01v8_lvt_GUWLND
X0 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X1 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X2 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X3 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X4 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X5 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X6 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X7 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
C0 out_left latch_right 0.1431f
C1 latch_left latch_right 5.15792f
C2 vinn tail 0.82695f
C3 vbias_p vinn 0.00222f
C4 vinn vout 0.12978f
C5 vbias_p tail 0.65167f
C6 tail vout 0.00803f
C7 vbias_p vout 0.14426f
C8 latch_right vinn 3.53507f
C9 latch_right tail 8.8942f
C10 vbias_p latch_right 0.00109f
C11 latch_right vout 0.72835f
C12 vdd vinp 4.26352f
C13 out_left vinp 0.22514f
C14 latch_left vinp 0.5043f
C15 out_left vdd 2.99708f
C16 vdd latch_left 1.3971f
C17 out_left latch_left 0.73463f
C18 vinn vinp 1.25697f
C19 tail vinp 2.91757f
C20 vbias_p vinp 0.03011f
C21 vout vinp 0.03655f
C22 vdd vinn 2.30474f
C23 vdd tail 2.22915f
C24 vbias_p vdd 2.11961f
C25 latch_right vinp 0.51311f
C26 vdd vout 1.62919f
C27 out_left vinn 0.08183f
C28 out_left tail 0.00652f
C29 out_left vbias_p 0.84152f
C30 out_left vout 0.6058f
C31 latch_left vinn 1.33911f
C32 latch_left tail 8.82993f
C33 vbias_p latch_left 0.00103f
C34 vdd latch_right 1.44611f
C35 latch_left vout 0.14014f
C36 vinp vss 0.4258f
C37 vinn vss 0.50566f
C38 tail vss 1.09774f
C39 vbias_p vss 0.82905f
C40 vdd vss 43.54159f
C41 vout vss 3.2381f
C42 latch_right vss 4.74799f
C43 out_left vss 3.38408f
C44 latch_left vss 5.11722f
.ends

.subckt sky130_fd_pr__pfet_01v8_A6MZLZ B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 G S 0.02934f
C1 D B 0.14266f
C2 D S 0.32105f
C3 B S 0.14266f
C4 G D 0.02934f
C5 G B 0.24043f
C6 S VSUBS 0.09023f
C7 D VSUBS 0.09023f
C8 G VSUBS 0.11914f
C9 B VSUBS 1.5811f
.ends

.subckt sky130_fd_pr__nfet_01v8_MH3LLV B D S G
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 S G 0.02545f
C1 D S 0.16211f
C2 D G 0.02545f
C3 S B 0.1317f
C4 D B 0.1317f
C5 G B 0.34289f
.ends

.subckt tmux_2to1 Y vdd XM5/G B A S vss
XXM1 vdd vdd XM5/G S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM2 vss vss XM5/G S sky130_fd_pr__nfet_01v8_MH3LLV
XXM3 vdd A Y S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM4 vss A Y XM5/G sky130_fd_pr__nfet_01v8_MH3LLV
XXM5 vdd Y B XM5/G vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM6 vss Y B S sky130_fd_pr__nfet_01v8_MH3LLV
C0 Y B 0.03022f
C1 vdd B 0.11322f
C2 A S 0.09932f
C3 XM5/G A 0.66126f
C4 Y vdd 0.18933f
C5 A Y 0.03022f
C6 A vdd 0.05809f
C7 XM5/G S 0.4752f
C8 S B 0.0426f
C9 XM5/G B 0.09611f
C10 Y S 0.13093f
C11 XM5/G Y 0.31571f
C12 vdd S 0.27839f
C13 XM5/G vdd 0.17343f
C14 B vss 0.39578f
C15 S vss 1.22376f
C16 Y vss 0.38976f
C17 XM5/G vss 0.68597f
C18 vdd vss 4.09633f
C19 A vss 0.18036f
.ends

.subckt sky130_fd_pr__res_generic_m1_SPQYYJ R1 R2 m1_n100_n100# VSUBS
R0 R1 R2 sky130_fd_pr__res_generic_m1 w=1 l=1
C0 R2 VSUBS 0.07104f
C1 R1 VSUBS 0.07104f
C2 m1_n100_n100# VSUBS 0.10692f
.ends

.subckt inv vin vdd vout vss
XXMn vss vss vout vin sky130_fd_pr__nfet_01v8_MH3LLV
XXMp vdd vdd vout vin vss sky130_fd_pr__pfet_01v8_A6MZLZ
C0 vin vout 0.12658f
C1 vdd vout 0.11998f
C2 vdd vin 0.13776f
C3 vin vss 0.56678f
C4 vout vss 0.40687f
C5 vdd vss 1.84972f
.ends

.subckt buffer in out vdd inv_1/vin vss
Xinv_0 in vdd inv_1/vin vss inv
Xinv_1 inv_1/vin vdd out vss inv
C0 vdd inv_1/vin 0.16476f
C1 out inv_1/vin 0.0071f
C2 out vdd 0.00589f
C3 in inv_1/vin 0.01628f
C4 vdd in 0.01965f
C5 inv_1/vin vss 0.60193f
C6 out vss 0.3255f
C7 in vss 0.41789f
C8 vdd vss 3.06334f
.ends

.subckt tmux_7therm_to_3bin d0 d1 d2 d3 d4 d5 d6 q0 q1 q2 buffer_7/inv_1/vin buffer_3/inv_1/vin
+ buffer_5/out buffer_2/out buffer_4/inv_1/vin buffer_0/inv_1/vin buffer_6/out R1/R2
+ buffer_0/out buffer_5/inv_1/vin buffer_1/inv_1/vin tmux_2to1_0/XM5/G R1/R1 tmux_2to1_3/A
+ tmux_2to1_3/XM5/G buffer_6/inv_1/vin buffer_2/inv_1/vin R1/m1_n100_n100# buffer_1/out
+ buffer_8/in vdd vss buffer_7/in buffer_4/out
Xtmux_2to1_1 buffer_8/in vdd tmux_2to1_1/XM5/G buffer_5/out buffer_1/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_2 tmux_2to1_3/B vdd tmux_2to1_2/XM5/G buffer_6/out buffer_2/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_3 buffer_7/in vdd tmux_2to1_3/XM5/G tmux_2to1_3/B tmux_2to1_3/A buffer_8/in
+ vss tmux_2to1
XR1 R1/R1 R1/R2 R1/m1_n100_n100# vss sky130_fd_pr__res_generic_m1_SPQYYJ
Xbuffer_0 d0 buffer_0/out vdd buffer_0/inv_1/vin vss buffer
Xbuffer_1 d1 buffer_1/out vdd buffer_1/inv_1/vin vss buffer
Xbuffer_2 d2 buffer_2/out vdd buffer_2/inv_1/vin vss buffer
Xbuffer_3 d3 R1/R2 vdd buffer_3/inv_1/vin vss buffer
Xbuffer_4 d4 buffer_4/out vdd buffer_4/inv_1/vin vss buffer
Xbuffer_5 d5 buffer_5/out vdd buffer_5/inv_1/vin vss buffer
Xbuffer_6 d6 buffer_6/out vdd buffer_6/inv_1/vin vss buffer
Xbuffer_7 buffer_7/in q0 vdd buffer_7/inv_1/vin vss buffer
Xbuffer_8 buffer_8/in q1 vdd buffer_8/inv_1/vin vss buffer
Xbuffer_9 R1/R1 q2 vdd buffer_9/inv_1/vin vss buffer
Xtmux_2to1_0 tmux_2to1_3/A vdd tmux_2to1_0/XM5/G buffer_4/out buffer_0/out R1/R1 vss
+ tmux_2to1
C0 tmux_2to1_3/XM5/G buffer_7/in 0.01403f
C1 tmux_2to1_3/B vdd 1.44834f
C2 buffer_4/out buffer_5/out 1.96436f
C3 vdd d3 0.07265f
C4 buffer_5/out buffer_1/out 0.05669f
C5 R1/R1 buffer_7/in 0.00295f
C6 buffer_6/out vdd 3.00774f
C7 tmux_2to1_3/B tmux_2to1_3/XM5/G 0.0457f
C8 d2 tmux_2to1_3/B 0
C9 buffer_0/inv_1/vin buffer_0/out 0.00873f
C10 d2 d3 0.00435f
C11 tmux_2to1_3/B R1/R1 0.24354f
C12 tmux_2to1_3/XM5/G vdd 0.0495f
C13 d3 R1/R1 0
C14 buffer_0/inv_1/vin buffer_1/inv_1/vin 0.00435f
C15 buffer_4/out buffer_7/in 0.04488f
C16 tmux_2to1_1/XM5/G buffer_5/out 0.02579f
C17 d2 vdd 0.07265f
C18 vdd d0 0.0683f
C19 tmux_2to1_0/XM5/G buffer_7/in 0.00597f
C20 buffer_6/out R1/R1 0.20693f
C21 d4 buffer_4/out 0.00133f
C22 buffer_1/out buffer_7/in 0
C23 d1 buffer_8/in 0
C24 d5 buffer_5/out 0.00133f
C25 vdd R1/R1 2.2016f
C26 buffer_2/out tmux_2to1_2/XM5/G 0.14365f
C27 tmux_2to1_3/B buffer_4/out 0.27941f
C28 buffer_5/inv_1/vin buffer_5/out 0.00827f
C29 buffer_2/inv_1/vin buffer_1/inv_1/vin 0.00438f
C30 buffer_8/inv_1/vin buffer_5/out 0
C31 tmux_2to1_3/B buffer_1/out 0
C32 tmux_2to1_3/B buffer_9/inv_1/vin 0.00176f
C33 tmux_2to1_3/XM5/G R1/R1 0
C34 d2 R1/R1 0.00119f
C35 buffer_6/out buffer_4/out 1.41966f
C36 buffer_4/inv_1/vin buffer_5/out 0
C37 d0 R1/R1 0
C38 tmux_2to1_3/A buffer_5/out 0.00456f
C39 buffer_4/out vdd 1.78677f
C40 buffer_8/in buffer_1/inv_1/vin 0
C41 R1/m1_n100_n100# buffer_5/out 0.01185f
C42 tmux_2to1_1/XM5/G buffer_7/in 0
C43 buffer_6/out buffer_9/inv_1/vin 0.00222f
C44 vdd tmux_2to1_0/XM5/G 0.05854f
C45 vdd buffer_1/out 0.83708f
C46 vdd buffer_9/inv_1/vin 0.03021f
C47 q1 buffer_7/in 0
C48 tmux_2to1_3/XM5/G buffer_4/out 0.04713f
C49 d4 d5 0.00435f
C50 tmux_2to1_1/XM5/G tmux_2to1_3/B 0
C51 tmux_2to1_3/XM5/G buffer_1/out 0
C52 buffer_8/inv_1/vin buffer_7/in 0
C53 q0 buffer_7/in 0
C54 R1/R2 buffer_5/out 0.01212f
C55 q1 tmux_2to1_3/B 0
C56 buffer_4/out R1/R1 0.26729f
C57 tmux_2to1_0/XM5/G d0 0
C58 tmux_2to1_3/A buffer_7/in 0.38438f
C59 tmux_2to1_0/XM5/G R1/R1 0.0674f
C60 buffer_1/out R1/R1 0.22519f
C61 buffer_3/inv_1/vin buffer_5/out 0
C62 tmux_2to1_1/XM5/G vdd 0.04059f
C63 buffer_9/inv_1/vin R1/R1 0.00349f
C64 buffer_8/inv_1/vin tmux_2to1_3/B 0.00974f
C65 d5 vdd 0.07265f
C66 q1 vdd 0.01294f
C67 buffer_6/out buffer_5/inv_1/vin 0
C68 tmux_2to1_3/A tmux_2to1_3/B 0.0101f
C69 buffer_5/inv_1/vin vdd 0.32846f
C70 buffer_8/in buffer_5/out 0.33947f
C71 buffer_8/inv_1/vin vdd 0.02538f
C72 buffer_4/out tmux_2to1_0/XM5/G 0.02654f
C73 vdd q0 0.01294f
C74 buffer_4/out buffer_1/out 0.00456f
C75 buffer_2/out buffer_5/out 0.05213f
C76 buffer_6/out buffer_4/inv_1/vin 0
C77 tmux_2to1_1/XM5/G R1/R1 0.13419f
C78 vdd buffer_4/inv_1/vin 0.32846f
C79 tmux_2to1_3/A vdd 0.31099f
C80 buffer_6/out R1/m1_n100_n100# 0
C81 R1/m1_n100_n100# vdd 0.01544f
C82 tmux_2to1_3/A tmux_2to1_3/XM5/G 0.04146f
C83 tmux_2to1_1/XM5/G buffer_4/out 0.02598f
C84 tmux_2to1_3/B buffer_2/inv_1/vin 0
C85 tmux_2to1_3/A d0 0
C86 buffer_0/inv_1/vin vdd 0.32203f
C87 buffer_8/in buffer_7/in 0.24628f
C88 buffer_6/out R1/R2 0.00154f
C89 tmux_2to1_1/XM5/G tmux_2to1_0/XM5/G 0.00433f
C90 tmux_2to1_3/A R1/R1 0.0222f
C91 R1/R2 vdd 0.32828f
C92 tmux_2to1_1/XM5/G buffer_1/out 0.18587f
C93 R1/m1_n100_n100# R1/R1 0.04565f
C94 buffer_6/out buffer_3/inv_1/vin 0
C95 tmux_2to1_2/XM5/G buffer_5/out 0.09828f
C96 buffer_3/inv_1/vin vdd 0.32836f
C97 q2 tmux_2to1_3/B 0
C98 buffer_6/out buffer_6/inv_1/vin 0.00786f
C99 buffer_2/inv_1/vin vdd 0.32649f
C100 tmux_2to1_3/B buffer_8/in 0.28179f
C101 vdd buffer_6/inv_1/vin 0.32835f
C102 buffer_2/out tmux_2to1_3/B 0.04026f
C103 buffer_0/inv_1/vin R1/R1 0.01886f
C104 buffer_4/out buffer_4/inv_1/vin 0.0079f
C105 tmux_2to1_3/A buffer_4/out 0.60354f
C106 buffer_8/inv_1/vin buffer_9/inv_1/vin 0.00438f
C107 R1/m1_n100_n100# buffer_4/out 0.00131f
C108 R1/R2 R1/R1 0.03366f
C109 q2 vdd 0.01294f
C110 tmux_2to1_3/A tmux_2to1_0/XM5/G 0.08101f
C111 buffer_6/out buffer_2/out 0.01539f
C112 vdd buffer_8/in 0.52301f
C113 tmux_2to1_3/A buffer_1/out 0
C114 buffer_2/out vdd 0.64599f
C115 buffer_3/inv_1/vin R1/R1 0.00894f
C116 buffer_2/inv_1/vin R1/R1 0.02182f
C117 tmux_2to1_3/XM5/G buffer_8/in 0.34642f
C118 buffer_0/out buffer_7/in 0
C119 R1/R2 buffer_4/out 0.00232f
C120 buffer_7/inv_1/vin buffer_7/in 0.00796f
C121 buffer_2/out d2 0
C122 buffer_0/inv_1/vin tmux_2to1_0/XM5/G 0
C123 q2 R1/R1 0
C124 tmux_2to1_3/B tmux_2to1_2/XM5/G 0.03416f
C125 buffer_8/in R1/R1 0.07792f
C126 tmux_2to1_3/A tmux_2to1_1/XM5/G 0
C127 buffer_3/inv_1/vin buffer_4/out 0
C128 buffer_2/out R1/R1 0.2789f
C129 buffer_6/out tmux_2to1_2/XM5/G 0.02333f
C130 d1 vdd 0.07265f
C131 buffer_5/inv_1/vin buffer_4/inv_1/vin 0.00435f
C132 vdd tmux_2to1_2/XM5/G 0.05427f
C133 tmux_2to1_3/A q0 0
C134 buffer_4/out buffer_8/in 0.18314f
C135 vdd buffer_0/out 0.83616f
C136 buffer_2/out buffer_4/out 0.0018f
C137 buffer_7/inv_1/vin vdd 0.02382f
C138 buffer_8/in buffer_1/out 0.06403f
C139 d2 d1 0.00438f
C140 d1 d0 0.00435f
C141 buffer_6/out d6 0.00132f
C142 d6 vdd 0.07265f
C143 vdd buffer_1/inv_1/vin 0.32649f
C144 d1 R1/R1 0
C145 tmux_2to1_2/XM5/G R1/R1 0.26532f
C146 buffer_0/out d0 0.0015f
C147 buffer_0/out R1/R1 0.11396f
C148 buffer_0/inv_1/vin tmux_2to1_3/A 0
C149 buffer_5/inv_1/vin buffer_6/inv_1/vin 0.00438f
C150 tmux_2to1_1/XM5/G buffer_8/in 0.12457f
C151 buffer_5/out buffer_7/in 0.00264f
C152 R1/m1_n100_n100# R1/R2 0.0386f
C153 buffer_3/inv_1/vin buffer_4/inv_1/vin 0.00438f
C154 buffer_4/out tmux_2to1_2/XM5/G 0.07683f
C155 buffer_1/inv_1/vin R1/R1 0.02062f
C156 q1 buffer_8/in 0
C157 R1/m1_n100_n100# buffer_3/inv_1/vin 0.00103f
C158 d1 buffer_1/out 0.00148f
C159 buffer_4/out buffer_0/out 0.0414f
C160 buffer_7/inv_1/vin buffer_4/out 0.00238f
C161 tmux_2to1_3/B buffer_5/out 0.16421f
C162 buffer_8/inv_1/vin buffer_8/in 0.01384f
C163 tmux_2to1_0/XM5/G buffer_0/out 0.18135f
C164 tmux_2to1_3/A buffer_8/in 0.1382f
C165 buffer_6/out buffer_5/out 0.48773f
C166 vdd buffer_5/out 1.96257f
C167 buffer_1/inv_1/vin buffer_1/out 0.0086f
C168 tmux_2to1_1/XM5/G tmux_2to1_2/XM5/G 0.00433f
C169 buffer_3/inv_1/vin buffer_2/inv_1/vin 0.00435f
C170 tmux_2to1_3/XM5/G buffer_5/out 0.01262f
C171 tmux_2to1_3/B buffer_7/in 0.20877f
C172 buffer_5/out R1/R1 0.55887f
C173 d4 d3 0.00438f
C174 vdd buffer_7/in 0.23539f
C175 buffer_2/out buffer_2/inv_1/vin 0.00356f
C176 d6 d5 0.00438f
C177 buffer_8/inv_1/vin buffer_7/inv_1/vin 0.00435f
C178 d4 vdd 0.07265f
C179 tmux_2to1_3/A buffer_0/out 0.05826f
C180 buffer_6/out tmux_2to1_3/B 0.18281f
C181 tmux_2to1_3/A buffer_7/inv_1/vin 0
C182 tmux_2to1_3/A vss 0.7137f
C183 tmux_2to1_0/XM5/G vss 0.55203f
C184 buffer_9/inv_1/vin vss 0.83718f
C185 q2 vss 0.40182f
C186 buffer_8/inv_1/vin vss 0.83586f
C187 q1 vss 0.40182f
C188 buffer_7/inv_1/vin vss 0.83588f
C189 q0 vss 0.40182f
C190 buffer_6/inv_1/vin vss 0.54713f
C191 buffer_6/out vss 1.08087f
C192 d6 vss 0.42023f
C193 buffer_5/inv_1/vin vss 0.54811f
C194 buffer_5/out vss 1.1426f
C195 d5 vss 0.41693f
C196 vdd vss 81.61826f
C197 buffer_4/inv_1/vin vss 0.54811f
C198 buffer_4/out vss 1.13891f
C199 d4 vss 0.41693f
C200 buffer_3/inv_1/vin vss 0.54811f
C201 R1/R2 vss 0.24595f
C202 d3 vss 0.41694f
C203 buffer_2/inv_1/vin vss 0.55981f
C204 buffer_2/out vss 0.38944f
C205 d2 vss 0.41693f
C206 buffer_1/inv_1/vin vss 0.55981f
C207 buffer_1/out vss 0.403f
C208 d1 vss 0.41693f
C209 buffer_0/inv_1/vin vss 0.55981f
C210 buffer_0/out vss 0.40723f
C211 d0 vss 0.42457f
C212 R1/m1_n100_n100# vss 0.11104f
C213 buffer_8/in vss 1.94693f
C214 buffer_7/in vss 1.30882f
C215 tmux_2to1_3/XM5/G vss 0.55181f
C216 R1/R1 vss 4.97016f
C217 tmux_2to1_3/B vss 1.00035f
C218 tmux_2to1_2/XM5/G vss 0.54992f
C219 tmux_2to1_1/XM5/G vss 0.55178f
.ends

.subckt flashADC_3bit_extracted vin vref dout0 dout1 dout2 d0 d1 d2 d3 d4 d5 d6 vdd
+ vss
Xvbias_generation_0 vbias_generation_0/bias_n vdd vbias_generation_0/XR_bias_2/R2
+ vbias_generation_0/XR_bias_4/R1 vbias_generation_0/XR_bias_3/R2 comp_p_6/vbias_p
+ vss vbias_generation
Xres_ladder_vref_0 comp_p_2/vinn comp_p_5/vinn comp_p_6/vinn vref comp_p_3/vinn comp_p_0/vinn
+ comp_p_1/vinn comp_p_4/vinn vss res_ladder_vref
Xcomp_p_1 vin comp_p_1/vinn comp_p_6/vbias_p vdd comp_p_1/tail d0 comp_p_1/latch_right
+ comp_p_1/out_left comp_p_1/latch_left vss comp_p
Xcomp_p_0 vin comp_p_0/vinn comp_p_6/vbias_p vdd comp_p_0/tail d1 comp_p_0/latch_right
+ comp_p_0/out_left comp_p_0/latch_left vss comp_p
Xcomp_p_2 vin comp_p_2/vinn comp_p_6/vbias_p vdd comp_p_2/tail d2 comp_p_2/latch_right
+ comp_p_2/out_left comp_p_2/latch_left vss comp_p
Xcomp_p_3 vin comp_p_3/vinn comp_p_6/vbias_p vdd comp_p_3/tail d3 comp_p_3/latch_right
+ comp_p_3/out_left comp_p_3/latch_left vss comp_p
Xcomp_p_4 vin comp_p_4/vinn comp_p_6/vbias_p vdd comp_p_4/tail d4 comp_p_4/latch_right
+ comp_p_4/out_left comp_p_4/latch_left vss comp_p
Xcomp_p_5 vin comp_p_5/vinn comp_p_6/vbias_p vdd comp_p_5/tail d5 comp_p_5/latch_right
+ comp_p_5/out_left comp_p_5/latch_left vss comp_p
Xcomp_p_6 vin comp_p_6/vinn comp_p_6/vbias_p vdd comp_p_6/tail d6 comp_p_6/latch_right
+ comp_p_6/out_left comp_p_6/latch_left vss comp_p
Xtmux_7therm_to_3bin_0 d0 d1 d2 d3 d4 d5 d6 dout0 dout1 dout2 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_3/inv_1/vin tmux_7therm_to_3bin_0/buffer_5/out tmux_7therm_to_3bin_0/buffer_2/out
+ tmux_7therm_to_3bin_0/buffer_4/inv_1/vin tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_6/out tmux_7therm_to_3bin_0/R1/R2 tmux_7therm_to_3bin_0/buffer_0/out
+ tmux_7therm_to_3bin_0/buffer_5/inv_1/vin tmux_7therm_to_3bin_0/buffer_1/inv_1/vin
+ tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G tmux_7therm_to_3bin_0/R1/R1 tmux_7therm_to_3bin_0/tmux_2to1_3/A
+ tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G tmux_7therm_to_3bin_0/buffer_6/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_2/inv_1/vin tmux_7therm_to_3bin_0/R1/m1_n100_n100#
+ tmux_7therm_to_3bin_0/buffer_1/out tmux_7therm_to_3bin_0/buffer_8/in vdd vss tmux_7therm_to_3bin_0/buffer_7/in
+ tmux_7therm_to_3bin_0/buffer_4/out tmux_7therm_to_3bin
X0 vdd comp_p_4/out_left.t2 d4 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X1 comp_p_4/out_left comp_p_4/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X2 vdd comp_p_6/out_left.t2 d6 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X3 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d1.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X4 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d6.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X5 comp_p_1/out_left comp_p_1/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X6 comp_p_2/tail vin.t10 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X7 comp_p_4/tail vin.t16 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X8 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d4.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X9 comp_p_2/tail vin.t9 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X10 vdd comp_p_6/vbias_p.t3 comp_p_0/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X11 comp_p_4/latch_left.t1 comp_p_4/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X12 comp_p_1/tail vin.t2 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X13 comp_p_3/latch_left comp_p_3/latch_right.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X14 comp_p_4/tail vin.t19 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X15 comp_p_5/latch_right comp_p_5/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X16 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d6.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X17 comp_p_2/latch_right comp_p_2/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X18 comp_p_2/tail vin.t11 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X19 vdd comp_p_6/vbias_p.t5 comp_p_3/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X20 comp_p_1/tail vin.t3 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X21 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d1.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X22 vdd comp_p_0/out_left.t0 comp_p_0/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X23 comp_p_2/latch_left.t1 comp_p_2/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X24 comp_p_3/out_left comp_p_3/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X25 vdd comp_p_6/vbias_p.t6 comp_p_4/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X26 comp_p_4/tail vin.t18 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X27 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin d3.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X28 comp_p_3/latch_left.t1 comp_p_3/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X29 vdd comp_p_6/vbias_p.t8 comp_p_6/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X30 comp_p_6/tail vin.t24 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X31 comp_p_0/tail vin.t6 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X32 vdd comp_p_6/out_left.t0 comp_p_6/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X33 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d2.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X34 comp_p_0/tail vin.t4 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X35 comp_p_3/tail vin.t12 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X36 vdd comp_p_4/out_left.t0 comp_p_4/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X37 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d2.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X38 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin d3.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X39 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d5.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X40 comp_p_0/tail vin.t7 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X41 comp_p_5/tail vin.t21 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X42 comp_p_6/latch_right comp_p_6/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X43 comp_p_1/latch_right comp_p_1/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X44 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d5.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X45 comp_p_0/tail vin.t5 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X46 comp_p_1/latch_left.t1 comp_p_1/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X47 vdd comp_p_6/vbias_p.t2 comp_p_1/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X48 vdd comp_p_0/out_left.t2 d1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X49 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d0.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X50 vdd comp_p_3/out_left.t2 d3 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X51 comp_p_4/latch_right comp_p_4/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X52 comp_p_5/out_left comp_p_5/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X53 vdd comp_p_6/vbias_p.t4 comp_p_2/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X54 comp_p_3/latch_right comp_p_3/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X55 comp_p_5/latch_left.t1 comp_p_5/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X56 comp_p_3/latch_right.t1 comp_p_3/latch_right.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X57 comp_p_6/tail vin.t25 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X58 comp_p_6/tail vin.t26 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X59 comp_p_2/tail vin.t8 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X60 comp_p_4/tail vin.t17 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X61 comp_p_5/tail vin.t20 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X62 comp_p_6/out_left comp_p_6/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X63 comp_p_3/tail vin.t13 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X64 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d0.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X65 d3 comp_p_3/latch_right.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X66 comp_p_3/tail vin.t14 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X67 vdd comp_p_6/vbias_p.t7 comp_p_5/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X68 comp_p_6/tail vin.t27 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X69 comp_p_2/out_left comp_p_2/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X70 vdd comp_p_3/out_left.t0 comp_p_3/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X71 comp_p_1/tail vin.t0 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X72 vdd comp_p_6/vbias_p.t0 comp_p_6/vbias_p.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X73 comp_p_5/tail vin.t23 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X74 comp_p_6/latch_left.t1 comp_p_6/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X75 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d4.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X76 comp_p_3/tail vin.t15 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X77 comp_p_5/tail vin.t22 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X78 comp_p_1/tail vin.t1 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
R0 comp_p_6/vbias_p.t0 comp_p_6/vbias_p.n6 337.106
R1 comp_p_6/vbias_p comp_p_6/vbias_p.t0 332.425
R2 comp_p_6/vbias_p comp_p_6/vbias_p.t2 178.793
R3 comp_p_6/vbias_p comp_p_6/vbias_p.t8 178.793
R4 comp_p_6/vbias_p.n2 comp_p_6/vbias_p.t7 172.639
R5 comp_p_6/vbias_p.n2 comp_p_6/vbias_p.t5 172.639
R6 comp_p_6/vbias_p.n3 comp_p_6/vbias_p.t6 172.639
R7 comp_p_6/vbias_p.n3 comp_p_6/vbias_p.t4 172.639
R8 comp_p_6/vbias_p.n0 comp_p_6/vbias_p.t3 172.639
R9 comp_p_6/vbias_p comp_p_6/vbias_p.t1 23.0294
R10 comp_p_6/vbias_p.n8 comp_p_6/vbias_p 8.71581
R11 comp_p_6/vbias_p.n0 comp_p_6/vbias_p 6.78896
R12 comp_p_6/vbias_p.n7 comp_p_6/vbias_p 4.65471
R13 comp_p_6/vbias_p.n1 comp_p_6/vbias_p 3.50247
R14 comp_p_6/vbias_p.n7 comp_p_6/vbias_p 3.11545
R15 comp_p_6/vbias_p comp_p_6/vbias_p.n8 2.28805
R16 comp_p_6/vbias_p.n5 comp_p_6/vbias_p.n1 2.21875
R17 comp_p_6/vbias_p comp_p_6/vbias_p.n5 2.14383
R18 comp_p_6/vbias_p.n1 comp_p_6/vbias_p.n0 2.08314
R19 comp_p_6/vbias_p.n3 comp_p_6/vbias_p 1.28874
R20 comp_p_6/vbias_p comp_p_6/vbias_p.n2 1.15992
R21 comp_p_6/vbias_p.n6 comp_p_6/vbias_p 0.802583
R22 comp_p_6/vbias_p.n4 comp_p_6/vbias_p 0.714721
R23 comp_p_6/vbias_p.n8 comp_p_6/vbias_p.n7 0.451639
R24 comp_p_6/vbias_p.n4 comp_p_6/vbias_p.n3 0.445699
R25 comp_p_6/vbias_p.n5 comp_p_6/vbias_p.n4 0.379389
R26 comp_p_6/vbias_p.n6 comp_p_6/vbias_p 0.0564593
R27 vss.n887 vss.n794 137199
R28 vss.n562 vss.n208 43219
R29 vss.n764 vss.n763 42544.4
R30 vss.n764 vss.n227 40078.3
R31 vss.n562 vss.n227 40078.3
R32 vss.n793 vss.n792 15045.2
R33 vss.n792 vss.n207 11496.8
R34 vss.n767 vss.n764 10982.3
R35 vss.n830 vss.n815 10261.4
R36 vss.n830 vss.n799 10261.4
R37 vss.n885 vss.n805 10261.4
R38 vss.n879 vss.n805 10261.4
R39 vss.n909 vss.n906 8494.18
R40 vss.n930 vss.n889 8494.18
R41 vss.n930 vss.n890 8494.18
R42 vss.n914 vss.n913 7120.97
R43 vss.n913 vss.n901 7120.97
R44 vss.n919 vss.n898 7120.97
R45 vss.n919 vss.n918 7120.97
R46 vss.n925 vss.n893 7120.97
R47 vss.n925 vss.n894 7120.97
R48 vss.n842 vss.n840 6385.12
R49 vss.n842 vss.n841 6385.12
R50 vss.n835 vss.n833 6385.12
R51 vss.n835 vss.n834 6385.12
R52 vss.n848 vss.n846 6385.12
R53 vss.n848 vss.n847 6385.12
R54 vss.n825 vss.n823 6385.12
R55 vss.n825 vss.n824 6385.12
R56 vss.n863 vss.n861 6385.12
R57 vss.n863 vss.n862 6385.12
R58 vss.n857 vss.n855 6385.12
R59 vss.n857 vss.n856 6385.12
R60 vss.n874 vss.n873 6385.12
R61 vss.n874 vss.n820 6385.12
R62 vss.n868 vss.n867 6385.12
R63 vss.n868 vss.n819 6385.12
R64 vss.n881 vss.n806 6385.12
R65 vss.n881 vss.n880 6385.12
R66 vss.n191 vss.n77 5440.68
R67 vss.n954 vss.n75 5440.68
R68 vss.n122 vss.n63 5440.68
R69 vss.n68 vss.n66 5440.68
R70 vss.n428 vss.n240 5440.68
R71 vss.n365 vss.n363 5440.68
R72 vss.n426 vss.n248 5440.68
R73 vss.n159 vss.n78 5255.26
R74 vss.n952 vss.n79 5255.26
R75 vss.n965 vss.n59 5255.26
R76 vss.n963 vss.n962 5255.26
R77 vss.n284 vss.n269 5255.26
R78 vss.n403 vss.n343 5255.26
R79 vss.n321 vss.n272 5255.26
R80 vss.n887 vss.n208 5235.57
R81 vss.n334 vss.n204 5116.21
R82 vss.n334 vss.n202 5116.21
R83 vss.n933 vss.n204 5116.21
R84 vss.n933 vss.n202 5116.21
R85 vss.n794 vss.n793 4892.83
R86 vss.n133 vss.n89 4536.79
R87 vss.n176 vss.n133 4536.79
R88 vss.n181 vss.n82 4536.79
R89 vss.n947 vss.n82 4536.79
R90 vss.n145 vss.n136 4536.79
R91 vss.n136 vss.n85 4536.79
R92 vss.n973 vss.n29 4536.79
R93 vss.n29 vss.n18 4536.79
R94 vss.n34 vss.n15 4536.79
R95 vss.n42 vss.n34 4536.79
R96 vss.n975 vss.n20 4536.79
R97 vss.n988 vss.n20 4536.79
R98 vss.n333 vss.n259 4536.79
R99 vss.n413 vss.n259 4536.79
R100 vss.n280 vss.n279 4536.79
R101 vss.n304 vss.n280 4536.79
R102 vss.n408 vss.n337 4536.79
R103 vss.n408 vss.n338 4536.79
R104 vss.n389 vss.n359 4536.79
R105 vss.n389 vss.n357 4536.79
R106 vss.n306 vss.n276 4536.79
R107 vss.n308 vss.n276 4536.79
R108 vss.n410 vss.n332 4536.79
R109 vss.n410 vss.n250 4536.79
R110 vss.n154 vss.n78 4131.21
R111 vss.n153 vss.n86 4131.21
R112 vss.n190 vss.n88 4131.21
R113 vss.n148 vss.n146 4131.21
R114 vss.n149 vss.n128 4131.21
R115 vss.n952 vss.n74 4131.21
R116 vss.n142 vss.n137 4131.21
R117 vss.n183 vss.n141 4131.21
R118 vss.n90 vss.n84 4131.21
R119 vss.n945 vss.n91 4131.21
R120 vss.n121 vss.n59 4131.21
R121 vss.n45 vss.n43 4131.21
R122 vss.n47 vss.n46 4131.21
R123 vss.n16 vss.n11 4131.21
R124 vss.n990 vss.n12 4131.21
R125 vss.n962 vss.n67 4131.21
R126 vss.n41 vss.n36 4131.21
R127 vss.n977 vss.n40 4131.21
R128 vss.n35 vss.n14 4131.21
R129 vss.n65 vss.n19 4131.21
R130 vss.n269 vss.n239 4131.21
R131 vss.n290 vss.n271 4131.21
R132 vss.n414 vss.n246 4131.21
R133 vss.n289 vss.n270 4131.21
R134 vss.n258 vss.n244 4131.21
R135 vss.n346 vss.n343 4131.21
R136 vss.n378 vss.n377 4131.21
R137 vss.n380 vss.n379 4131.21
R138 vss.n352 vss.n345 4131.21
R139 vss.n386 vss.n366 4131.21
R140 vss.n321 vss.n247 4131.21
R141 vss.n323 vss.n266 4131.21
R142 vss.n262 vss.n242 4131.21
R143 vss.n316 vss.n268 4131.21
R144 vss.n327 vss.n243 4131.21
R145 vss.n694 vss.n693 4116.13
R146 vss.n154 vss.n77 3945.79
R147 vss.n158 vss.n86 3945.79
R148 vss.n153 vss.n88 3945.79
R149 vss.n150 vss.n146 3945.79
R150 vss.n149 vss.n148 3945.79
R151 vss.n954 vss.n74 3945.79
R152 vss.n177 vss.n142 3945.79
R153 vss.n183 vss.n137 3945.79
R154 vss.n84 vss.n83 3945.79
R155 vss.n945 vss.n90 3945.79
R156 vss.n122 vss.n121 3945.79
R157 vss.n48 vss.n43 3945.79
R158 vss.n47 vss.n45 3945.79
R159 vss.n60 vss.n16 3945.79
R160 vss.n990 vss.n11 3945.79
R161 vss.n68 vss.n67 3945.79
R162 vss.n41 vss.n26 3945.79
R163 vss.n977 vss.n36 3945.79
R164 vss.n21 vss.n14 3945.79
R165 vss.n35 vss.n19 3945.79
R166 vss.n428 vss.n239 3945.79
R167 vss.n297 vss.n271 3945.79
R168 vss.n290 vss.n246 3945.79
R169 vss.n281 vss.n270 3945.79
R170 vss.n289 vss.n244 3945.79
R171 vss.n363 vss.n346 3945.79
R172 vss.n377 vss.n370 3945.79
R173 vss.n380 vss.n378 3945.79
R174 vss.n352 vss.n342 3945.79
R175 vss.n386 vss.n345 3945.79
R176 vss.n426 vss.n247 3945.79
R177 vss.n323 vss.n265 3945.79
R178 vss.n266 vss.n242 3945.79
R179 vss.n278 vss.n268 3945.79
R180 vss.n316 vss.n243 3945.79
R181 vss.n820 vss.n812 3876.26
R182 vss.n862 vss.n812 3876.26
R183 vss.n847 vss.n814 3876.26
R184 vss.n841 vss.n814 3876.26
R185 vss.n834 vss.n815 3876.26
R186 vss.n840 vss.n801 3876.26
R187 vss.n833 vss.n801 3876.26
R188 vss.n833 vss.n799 3876.26
R189 vss.n841 vss.n816 3876.26
R190 vss.n834 vss.n816 3876.26
R191 vss.n823 vss.n802 3876.26
R192 vss.n846 vss.n802 3876.26
R193 vss.n846 vss.n798 3876.26
R194 vss.n840 vss.n798 3876.26
R195 vss.n856 vss.n813 3876.26
R196 vss.n824 vss.n813 3876.26
R197 vss.n824 vss.n817 3876.26
R198 vss.n847 vss.n817 3876.26
R199 vss.n861 vss.n803 3876.26
R200 vss.n855 vss.n803 3876.26
R201 vss.n855 vss.n797 3876.26
R202 vss.n823 vss.n797 3876.26
R203 vss.n862 vss.n818 3876.26
R204 vss.n856 vss.n818 3876.26
R205 vss.n867 vss.n804 3876.26
R206 vss.n873 vss.n804 3876.26
R207 vss.n873 vss.n796 3876.26
R208 vss.n861 vss.n796 3876.26
R209 vss.n880 vss.n810 3876.26
R210 vss.n819 vss.n810 3876.26
R211 vss.n877 vss.n819 3876.26
R212 vss.n877 vss.n820 3876.26
R213 vss.n885 vss.n806 3876.26
R214 vss.n806 vss.n795 3876.26
R215 vss.n867 vss.n795 3876.26
R216 vss.n880 vss.n879 3876.26
R217 vss.n158 vss.n89 3227.32
R218 vss.n176 vss.n150 3227.32
R219 vss.n147 vss.n128 3227.32
R220 vss.n181 vss.n177 3227.32
R221 vss.n145 vss.n141 3227.32
R222 vss.n947 vss.n83 3227.32
R223 vss.n91 vss.n85 3227.32
R224 vss.n973 vss.n48 3227.32
R225 vss.n46 vss.n44 3227.32
R226 vss.n60 vss.n18 3227.32
R227 vss.n975 vss.n26 3227.32
R228 vss.n42 vss.n40 3227.32
R229 vss.n988 vss.n21 3227.32
R230 vss.n65 vss.n15 3227.32
R231 vss.n297 vss.n279 3227.32
R232 vss.n414 vss.n413 3227.32
R233 vss.n304 vss.n281 3227.32
R234 vss.n333 vss.n258 3227.32
R235 vss.n370 vss.n337 3227.32
R236 vss.n379 vss.n359 3227.32
R237 vss.n342 vss.n338 3227.32
R238 vss.n366 vss.n357 3227.32
R239 vss.n306 vss.n265 3227.32
R240 vss.n332 vss.n262 3227.32
R241 vss.n308 vss.n278 3227.32
R242 vss.n327 vss.n250 3227.32
R243 vss.n495 vss.n208 2684.15
R244 vss.n887 vss.n207 2649.46
R245 vss.n503 vss.n485 2306.06
R246 vss.n494 vss.n485 2306.06
R247 vss.n503 vss.n486 2306.06
R248 vss.n494 vss.n486 2306.06
R249 vss.n513 vss.n475 2306.06
R250 vss.n505 vss.n475 2306.06
R251 vss.n513 vss.n476 2306.06
R252 vss.n505 vss.n476 2306.06
R253 vss.n616 vss.n612 2306.06
R254 vss.n616 vss.n613 2306.06
R255 vss.n626 vss.n470 2306.06
R256 vss.n471 vss.n470 2306.06
R257 vss.n578 vss.n550 2306.06
R258 vss.n593 vss.n550 2306.06
R259 vss.n578 vss.n551 2306.06
R260 vss.n593 vss.n551 2306.06
R261 vss.n564 vss.n557 2306.06
R262 vss.n575 vss.n557 2306.06
R263 vss.n564 vss.n558 2306.06
R264 vss.n575 vss.n558 2306.06
R265 vss.n492 vss.n483 2306.06
R266 vss.n496 vss.n492 2306.06
R267 vss.n493 vss.n483 2306.06
R268 vss.n496 vss.n493 2306.06
R269 vss.n481 vss.n473 2306.06
R270 vss.n507 vss.n481 2306.06
R271 vss.n482 vss.n473 2306.06
R272 vss.n507 vss.n482 2306.06
R273 vss.n618 vss.n528 2306.06
R274 vss.n618 vss.n532 2306.06
R275 vss.n624 vss.n517 2306.06
R276 vss.n517 vss.n472 2306.06
R277 vss.n590 vss.n586 2306.06
R278 vss.n590 vss.n587 2306.06
R279 vss.n609 vss.n534 2306.06
R280 vss.n609 vss.n535 2306.06
R281 vss.n580 vss.n553 2306.06
R282 vss.n584 vss.n553 2306.06
R283 vss.n580 vss.n554 2306.06
R284 vss.n584 vss.n554 2306.06
R285 vss.n566 vss.n561 2306.06
R286 vss.n561 vss.n556 2306.06
R287 vss.n567 vss.n566 2306.06
R288 vss.n567 vss.n556 2306.06
R289 vss.n740 vss.n720 2306.06
R290 vss.n729 vss.n720 2306.06
R291 vss.n740 vss.n721 2306.06
R292 vss.n729 vss.n721 2306.06
R293 vss.n711 vss.n646 2306.06
R294 vss.n743 vss.n646 2306.06
R295 vss.n711 vss.n647 2306.06
R296 vss.n743 vss.n647 2306.06
R297 vss.n698 vss.n667 2306.06
R298 vss.n696 vss.n667 2306.06
R299 vss.n708 vss.n652 2306.06
R300 vss.n708 vss.n653 2306.06
R301 vss.n680 vss.n669 2306.06
R302 vss.n692 vss.n669 2306.06
R303 vss.n680 vss.n670 2306.06
R304 vss.n692 vss.n670 2306.06
R305 vss.n676 vss.n673 2306.06
R306 vss.n683 vss.n673 2306.06
R307 vss.n676 vss.n674 2306.06
R308 vss.n683 vss.n674 2306.06
R309 vss.n727 vss.n718 2306.06
R310 vss.n731 vss.n727 2306.06
R311 vss.n728 vss.n718 2306.06
R312 vss.n731 vss.n728 2306.06
R313 vss.n713 vss.n649 2306.06
R314 vss.n717 vss.n649 2306.06
R315 vss.n713 vss.n650 2306.06
R316 vss.n717 vss.n650 2306.06
R317 vss.n440 vss.n438 2306.06
R318 vss.n446 vss.n438 2306.06
R319 vss.n445 vss.n440 2306.06
R320 vss.n446 vss.n445 2306.06
R321 vss.n762 vss.n229 2306.06
R322 vss.n441 vss.n229 2306.06
R323 vss.n762 vss.n230 2306.06
R324 vss.n441 vss.n230 2306.06
R325 vss.n779 vss.n213 2306.06
R326 vss.n790 vss.n213 2306.06
R327 vss.n779 vss.n214 2306.06
R328 vss.n790 vss.n214 2306.06
R329 vss.n766 vss.n220 2306.06
R330 vss.n776 vss.n220 2306.06
R331 vss.n766 vss.n221 2306.06
R332 vss.n776 vss.n221 2306.06
R333 vss.n781 vss.n217 2306.06
R334 vss.n217 vss.n212 2306.06
R335 vss.n782 vss.n781 2306.06
R336 vss.n782 vss.n212 2306.06
R337 vss.n768 vss.n226 2306.06
R338 vss.n226 vss.n219 2306.06
R339 vss.n769 vss.n768 2306.06
R340 vss.n769 vss.n219 2306.06
R341 vss.n888 vss.n206 2024.56
R342 vss.n190 vss.n87 1825.15
R343 vss.n117 vss.n12 1825.15
R344 vss.n322 vss.n241 1455.1
R345 vss.n427 vss.n245 1455.1
R346 vss.n467 vss.n463 1390.59
R347 vss.n467 vss.n457 1390.59
R348 vss.n464 vss.n462 1390.59
R349 vss.n464 vss.n456 1390.59
R350 vss.n520 vss.n516 1390.59
R351 vss.n520 vss.n519 1390.59
R352 vss.n530 vss.n529 1390.59
R353 vss.n531 vss.n530 1390.59
R354 vss.n544 vss.n543 1390.59
R355 vss.n543 vss.n539 1390.59
R356 vss.n545 vss.n542 1390.59
R357 vss.n545 vss.n538 1390.59
R358 vss.n663 vss.n662 1390.59
R359 vss.n662 vss.n658 1390.59
R360 vss.n664 vss.n661 1390.59
R361 vss.n664 vss.n657 1390.59
R362 vss.n322 vss.n267 1389.8
R363 vss.n427 vss.n241 1389.8
R364 vss.n914 vss.n903 1373.21
R365 vss.n918 vss.n917 1373.21
R366 vss.n917 vss.n901 1373.21
R367 vss.n909 vss.n901 1373.21
R368 vss.n922 vss.n893 1373.21
R369 vss.n922 vss.n898 1373.21
R370 vss.n915 vss.n898 1373.21
R371 vss.n915 vss.n914 1373.21
R372 vss.n893 vss.n889 1373.21
R373 vss.n894 vss.n890 1373.21
R374 vss.n896 vss.n894 1373.21
R375 vss.n918 vss.n896 1373.21
R376 vss.n150 vss.n135 1309.47
R377 vss.n158 vss.n135 1309.47
R378 vss.n148 vss.n134 1309.47
R379 vss.n153 vss.n134 1309.47
R380 vss.n159 vss.n158 1309.47
R381 vss.n155 vss.n153 1309.47
R382 vss.n155 vss.n154 1309.47
R383 vss.n189 vss.n128 1309.47
R384 vss.n190 vss.n189 1309.47
R385 vss.n191 vss.n190 1309.47
R386 vss.n83 vss.n79 1309.47
R387 vss.n92 vss.n90 1309.47
R388 vss.n92 vss.n74 1309.47
R389 vss.n91 vss.n75 1309.47
R390 vss.n141 vss.n132 1309.47
R391 vss.n132 vss.n91 1309.47
R392 vss.n187 vss.n137 1309.47
R393 vss.n187 vss.n90 1309.47
R394 vss.n177 vss.n131 1309.47
R395 vss.n131 vss.n83 1309.47
R396 vss.n121 vss.n64 1309.47
R397 vss.n64 vss.n11 1309.47
R398 vss.n965 vss.n60 1309.47
R399 vss.n63 vss.n12 1309.47
R400 vss.n60 vss.n33 1309.47
R401 vss.n48 vss.n33 1309.47
R402 vss.n30 vss.n11 1309.47
R403 vss.n45 vss.n30 1309.47
R404 vss.n32 vss.n12 1309.47
R405 vss.n46 vss.n32 1309.47
R406 vss.n67 vss.n62 1309.47
R407 vss.n62 vss.n35 1309.47
R408 vss.n963 vss.n21 1309.47
R409 vss.n66 vss.n65 1309.47
R410 vss.n983 vss.n21 1309.47
R411 vss.n983 vss.n26 1309.47
R412 vss.n981 vss.n35 1309.47
R413 vss.n981 vss.n36 1309.47
R414 vss.n65 vss.n28 1309.47
R415 vss.n40 vss.n28 1309.47
R416 vss.n328 vss.n262 1309.47
R417 vss.n328 vss.n327 1309.47
R418 vss.n288 vss.n239 1309.47
R419 vss.n289 vss.n288 1309.47
R420 vss.n284 vss.n281 1309.47
R421 vss.n258 vss.n240 1309.47
R422 vss.n298 vss.n281 1309.47
R423 vss.n298 vss.n297 1309.47
R424 vss.n291 vss.n289 1309.47
R425 vss.n291 vss.n290 1309.47
R426 vss.n415 vss.n258 1309.47
R427 vss.n415 vss.n414 1309.47
R428 vss.n403 vss.n342 1309.47
R429 vss.n400 vss.n345 1309.47
R430 vss.n400 vss.n346 1309.47
R431 vss.n366 vss.n365 1309.47
R432 vss.n379 vss.n361 1309.47
R433 vss.n366 vss.n361 1309.47
R434 vss.n378 vss.n369 1309.47
R435 vss.n369 vss.n345 1309.47
R436 vss.n374 vss.n370 1309.47
R437 vss.n374 vss.n342 1309.47
R438 vss.n278 vss.n272 1309.47
R439 vss.n317 vss.n316 1309.47
R440 vss.n317 vss.n247 1309.47
R441 vss.n327 vss.n248 1309.47
R442 vss.n315 vss.n266 1309.47
R443 vss.n316 vss.n315 1309.47
R444 vss.n277 vss.n265 1309.47
R445 vss.n278 vss.n277 1309.47
R446 vss.n117 vss.n116 1251.53
R447 vss.n307 vss.n210 1136.73
R448 vss.n307 vss.n267 1136.73
R449 vss.n412 vss.n245 1136.73
R450 vss.n412 vss.n411 1136.73
R451 vss.n888 vss.n887 1030.43
R452 vss.n612 vss.n462 915.471
R453 vss.n630 vss.n462 915.471
R454 vss.n630 vss.n463 915.471
R455 vss.n626 vss.n463 915.471
R456 vss.n613 vss.n456 915.471
R457 vss.n632 vss.n456 915.471
R458 vss.n632 vss.n457 915.471
R459 vss.n471 vss.n457 915.471
R460 vss.n529 vss.n528 915.471
R461 vss.n529 vss.n461 915.471
R462 vss.n516 vss.n461 915.471
R463 vss.n624 vss.n516 915.471
R464 vss.n532 vss.n531 915.471
R465 vss.n531 vss.n459 915.471
R466 vss.n519 vss.n459 915.471
R467 vss.n519 vss.n472 915.471
R468 vss.n586 vss.n542 915.471
R469 vss.n602 vss.n542 915.471
R470 vss.n602 vss.n544 915.471
R471 vss.n544 vss.n534 915.471
R472 vss.n587 vss.n538 915.471
R473 vss.n604 vss.n538 915.471
R474 vss.n604 vss.n539 915.471
R475 vss.n539 vss.n535 915.471
R476 vss.n698 vss.n661 915.471
R477 vss.n703 vss.n661 915.471
R478 vss.n703 vss.n663 915.471
R479 vss.n663 vss.n652 915.471
R480 vss.n696 vss.n657 915.471
R481 vss.n705 vss.n657 915.471
R482 vss.n705 vss.n658 915.471
R483 vss.n658 vss.n653 915.471
R484 vss.n411 vss.n409 751.02
R485 vss.n936 vss.n935 705.364
R486 vss.n831 vss.n829 666.73
R487 vss vss.n831 666.73
R488 vss.n409 vss.n336 659.184
R489 vss.n884 vss.n807 621.553
R490 vss vss.n811 619.196
R491 vss.n935 vss.n934 599.019
R492 vss.n116 vss.n5 585
R493 vss.n116 vss.n17 585
R494 vss.n118 vss.n117 585
R495 vss.n117 vss.n13 585
R496 vss.n767 vss.n218 560.645
R497 vss.n777 vss.n218 560.645
R498 vss.n780 vss.n211 560.645
R499 vss.n791 vss.n211 560.645
R500 vss.n678 vss.n677 560.645
R501 vss.n682 vss.n678 560.645
R502 vss.n681 vss.n668 560.645
R503 vss.n693 vss.n668 560.645
R504 vss.n697 vss.n694 560.645
R505 vss.n697 vss.n659 560.645
R506 vss.n704 vss.n659 560.645
R507 vss.n704 vss.n660 560.645
R508 vss.n660 vss.n651 560.645
R509 vss.n709 vss.n651 560.645
R510 vss.n712 vss.n648 560.645
R511 vss.n742 vss.n648 560.645
R512 vss.n741 vss.n719 560.645
R513 vss.n730 vss.n719 560.645
R514 vss.n565 vss.n555 560.645
R515 vss.n576 vss.n555 560.645
R516 vss.n579 vss.n552 560.645
R517 vss.n592 vss.n552 560.645
R518 vss.n591 vss.n585 560.645
R519 vss.n585 vss.n540 560.645
R520 vss.n603 vss.n540 560.645
R521 vss.n603 vss.n541 560.645
R522 vss.n541 vss.n533 560.645
R523 vss.n610 vss.n533 560.645
R524 vss.n617 vss.n611 560.645
R525 vss.n611 vss.n458 560.645
R526 vss.n631 vss.n458 560.645
R527 vss.n631 vss.n460 560.645
R528 vss.n625 vss.n460 560.645
R529 vss.n625 vss.n515 560.645
R530 vss.n514 vss.n474 560.645
R531 vss.n506 vss.n474 560.645
R532 vss.n504 vss.n484 560.645
R533 vss.n495 vss.n484 560.645
R534 vss.n905 vss 551.907
R535 vss.n910 vss.n905 551.907
R536 vss.n929 vss.n928 551.907
R537 vss.n336 vss.n335 550.859
R538 vss.n52 vss.n31 534.431
R539 vss.n169 vss.n130 531.552
R540 vss.n677 vss.n227 514.516
R541 vss.n565 vss.n562 514.516
R542 vss.n388 vss.n360 490.01
R543 vss.n388 vss.n387 490.01
R544 vss.n387 vss.n362 490.01
R545 vss.n362 vss.n206 490.01
R546 vss.n912 vss.n904 462.683
R547 vss.n912 vss.n911 462.683
R548 vss.n921 vss.n920 462.683
R549 vss.n920 vss.n900 462.683
R550 vss.n926 vss.n892 462.683
R551 vss.n927 vss.n926 462.683
R552 vss.n924 vss.n895 435.882
R553 vss.n924 vss.n923 435.882
R554 vss.n923 vss.n897 435.882
R555 vss.n916 vss.n897 435.882
R556 vss.n916 vss.n902 435.882
R557 vss.n908 vss.n902 435.882
R558 vss.n907 vss.n906 424.591
R559 vss.n376 vss.n375 417.005
R560 vss.n375 vss.n344 417.005
R561 vss.n402 vss.n344 417.005
R562 vss.n402 vss.n401 417.005
R563 vss.n335 vss.n205 417.005
R564 vss.n932 vss.n205 417.005
R565 vss.n837 vss.n836 414.872
R566 vss.n836 vss.n832 414.872
R567 vss.n843 vss.n839 414.872
R568 vss.n844 vss.n843 414.872
R569 vss.n852 vss.n826 414.872
R570 vss.n828 vss.n826 414.872
R571 vss.n850 vss.n849 414.872
R572 vss.n849 vss.n845 414.872
R573 vss.n858 vss.n854 414.872
R574 vss.n859 vss.n858 414.872
R575 vss.n865 vss.n864 414.872
R576 vss.n864 vss.n860 414.872
R577 vss.n870 vss.n869 414.872
R578 vss.n869 vss.n821 414.872
R579 vss.n875 vss.n872 414.872
R580 vss.n876 vss.n875 414.872
R581 vss.n883 vss.n882 414.872
R582 vss.n882 vss.n809 414.872
R583 vss.n712 vss.n709 376.13
R584 vss.n592 vss.n591 376.13
R585 vss.n617 vss.n610 376.13
R586 vss.n515 vss.n514 376.13
R587 vss.n780 vss.n777 369.033
R588 vss.n682 vss.n681 369.033
R589 vss.n742 vss.n741 369.033
R590 vss.n579 vss.n576 369.033
R591 vss.n506 vss.n504 369.033
R592 vss.n620 vss.n619 343.154
R593 vss.n895 vss.n888 339.783
R594 vss vss.n203 335.06
R595 vss.n886 vss.n800 302.937
R596 vss.n878 vss.n800 302.937
R597 vss.n331 vss.n251 294.776
R598 vss.n286 vss.n282 294.776
R599 vss.n261 vss.n260 294.776
R600 vss.n972 vss.n49 294.776
R601 vss.n175 vss.n151 294.776
R602 vss.n144 vss.n143 294.776
R603 vss.n974 vss.n22 294.776
R604 vss.n111 vss.n110 294.776
R605 vss.n180 vss.n81 294.776
R606 vss.n390 vss.n358 294.776
R607 vss.n407 vss.n339 294.776
R608 vss.n305 vss.n275 294.776
R609 vss.n770 vss.n769 292.5
R610 vss.n769 vss.n218 292.5
R611 vss.n226 vss 292.5
R612 vss.n226 vss.n218 292.5
R613 vss.n783 vss.n782 292.5
R614 vss.n782 vss.n211 292.5
R615 vss.n217 vss 292.5
R616 vss.n217 vss.n211 292.5
R617 vss vss.n221 292.5
R618 vss.n221 vss.n218 292.5
R619 vss.n222 vss.n220 292.5
R620 vss.n220 vss.n218 292.5
R621 vss vss.n214 292.5
R622 vss.n214 vss.n211 292.5
R623 vss.n215 vss.n213 292.5
R624 vss.n213 vss.n211 292.5
R625 vss vss.n230 292.5
R626 vss.n230 vss.n228 292.5
R627 vss.n231 vss.n229 292.5
R628 vss.n229 vss.n228 292.5
R629 vss.n445 vss 292.5
R630 vss.n445 vss.n444 292.5
R631 vss.n438 vss.n437 292.5
R632 vss.n444 vss.n438 292.5
R633 vss.n715 vss.n650 292.5
R634 vss.n650 vss.n648 292.5
R635 vss vss.n649 292.5
R636 vss.n649 vss.n648 292.5
R637 vss.n728 vss.n726 292.5
R638 vss.n728 vss.n719 292.5
R639 vss.n727 vss 292.5
R640 vss.n727 vss.n719 292.5
R641 vss.n674 vss 292.5
R642 vss.n678 vss.n674 292.5
R643 vss.n673 vss.n672 292.5
R644 vss.n678 vss.n673 292.5
R645 vss vss.n670 292.5
R646 vss.n670 vss.n668 292.5
R647 vss.n671 vss.n669 292.5
R648 vss.n669 vss.n668 292.5
R649 vss vss.n653 292.5
R650 vss.n653 vss.n651 292.5
R651 vss vss.n705 292.5
R652 vss.n705 vss.n704 292.5
R653 vss.n696 vss 292.5
R654 vss.n697 vss.n696 292.5
R655 vss.n699 vss.n698 292.5
R656 vss.n698 vss.n697 292.5
R657 vss.n703 vss.n702 292.5
R658 vss.n704 vss.n703 292.5
R659 vss.n654 vss.n652 292.5
R660 vss.n652 vss.n651 292.5
R661 vss.n647 vss 292.5
R662 vss.n648 vss.n647 292.5
R663 vss.n646 vss.n645 292.5
R664 vss.n648 vss.n646 292.5
R665 vss vss.n721 292.5
R666 vss.n721 vss.n719 292.5
R667 vss.n722 vss.n720 292.5
R668 vss.n720 vss.n719 292.5
R669 vss.n568 vss.n567 292.5
R670 vss.n567 vss.n555 292.5
R671 vss.n561 vss 292.5
R672 vss.n561 vss.n555 292.5
R673 vss.n582 vss.n554 292.5
R674 vss.n554 vss.n552 292.5
R675 vss vss.n553 292.5
R676 vss.n553 vss.n552 292.5
R677 vss.n607 vss.n535 292.5
R678 vss.n535 vss.n533 292.5
R679 vss.n605 vss.n604 292.5
R680 vss.n604 vss.n603 292.5
R681 vss.n588 vss.n587 292.5
R682 vss.n587 vss.n585 292.5
R683 vss vss.n586 292.5
R684 vss.n586 vss.n585 292.5
R685 vss.n602 vss 292.5
R686 vss.n603 vss.n602 292.5
R687 vss vss.n534 292.5
R688 vss.n534 vss.n533 292.5
R689 vss.n523 vss.n472 292.5
R690 vss.n625 vss.n472 292.5
R691 vss.n525 vss.n459 292.5
R692 vss.n631 vss.n459 292.5
R693 vss.n532 vss.n527 292.5
R694 vss.n611 vss.n532 292.5
R695 vss.n528 vss 292.5
R696 vss.n611 vss.n528 292.5
R697 vss vss.n461 292.5
R698 vss.n631 vss.n461 292.5
R699 vss.n624 vss 292.5
R700 vss.n625 vss.n624 292.5
R701 vss.n482 vss.n480 292.5
R702 vss.n482 vss.n474 292.5
R703 vss.n481 vss 292.5
R704 vss.n481 vss.n474 292.5
R705 vss.n493 vss.n491 292.5
R706 vss.n493 vss.n484 292.5
R707 vss.n492 vss 292.5
R708 vss.n492 vss.n484 292.5
R709 vss vss.n558 292.5
R710 vss.n558 vss.n555 292.5
R711 vss.n559 vss.n557 292.5
R712 vss.n557 vss.n555 292.5
R713 vss.n551 vss 292.5
R714 vss.n552 vss.n551 292.5
R715 vss.n550 vss.n549 292.5
R716 vss.n552 vss.n550 292.5
R717 vss.n471 vss 292.5
R718 vss.n625 vss.n471 292.5
R719 vss vss.n632 292.5
R720 vss.n632 vss.n631 292.5
R721 vss vss.n613 292.5
R722 vss.n613 vss.n611 292.5
R723 vss.n614 vss.n612 292.5
R724 vss.n612 vss.n611 292.5
R725 vss.n630 vss.n629 292.5
R726 vss.n631 vss.n630 292.5
R727 vss.n627 vss.n626 292.5
R728 vss.n626 vss.n625 292.5
R729 vss vss.n476 292.5
R730 vss.n476 vss.n474 292.5
R731 vss.n477 vss.n475 292.5
R732 vss.n475 vss.n474 292.5
R733 vss vss.n486 292.5
R734 vss.n486 vss.n484 292.5
R735 vss.n487 vss.n485 292.5
R736 vss.n485 vss.n484 292.5
R737 vss vss.n201 285.604
R738 vss.n429 vss.n238 280.32
R739 vss.n123 vss.n120 280.32
R740 vss.n193 vss.n192 280.32
R741 vss.n105 vss.n69 280.32
R742 vss.n955 vss.n73 280.32
R743 vss.n364 vss.n348 280.32
R744 vss.n425 vss.n424 280.32
R745 vss.n283 vss.n237 268.425
R746 vss.n295 vss.n294 268.425
R747 vss.n293 vss.n257 268.425
R748 vss.n56 vss.n55 268.425
R749 vss.n54 vss.n53 268.425
R750 vss.n115 vss.n58 268.425
R751 vss.n157 vss.n126 268.425
R752 vss.n173 vss.n172 268.425
R753 vss.n171 vss.n170 268.425
R754 vss.n979 vss.n38 268.425
R755 vss.n978 vss.n39 268.425
R756 vss.n961 vss.n960 268.425
R757 vss.n951 vss.n72 268.425
R758 vss.n185 vss.n138 268.425
R759 vss.n184 vss.n140 268.425
R760 vss.n398 vss.n341 268.425
R761 vss.n371 vss.n367 268.425
R762 vss.n382 vss.n381 268.425
R763 vss.n320 vss.n319 268.425
R764 vss.n325 vss.n324 268.425
R765 vss.n330 vss.n326 268.425
R766 vss.n285 vss.n283 268.274
R767 vss.n966 vss.n58 268.274
R768 vss.n160 vss.n157 268.274
R769 vss.n961 vss.n23 268.274
R770 vss.n951 vss.n950 268.274
R771 vss.n404 vss.n341 268.274
R772 vss.n320 vss.n273 268.274
R773 vss.n296 vss.n295 256.377
R774 vss.n294 vss.n293 256.377
R775 vss.n971 vss.n56 256.377
R776 vss.n55 vss.n54 256.377
R777 vss.n174 vss.n173 256.377
R778 vss.n172 vss.n171 256.377
R779 vss.n38 vss.n25 256.377
R780 vss.n979 vss.n978 256.377
R781 vss.n179 vss.n138 256.377
R782 vss.n185 vss.n184 256.377
R783 vss.n372 vss.n371 256.377
R784 vss.n381 vss.n367 256.377
R785 vss.n324 vss.n264 256.377
R786 vss.n326 vss.n325 256.377
R787 vss.n430 vss.n429 256
R788 vss.n124 vss.n123 256
R789 vss.n194 vss.n193 256
R790 vss.n958 vss.n69 256
R791 vss.n956 vss.n955 256
R792 vss.n397 vss.n348 256
R793 vss.n425 vss.n235 256
R794 vss.n883 vss.n808 251.859
R795 vss.n870 vss.n808 251.859
R796 vss.n854 vss.n853 251.859
R797 vss.n853 vss.n852 251.859
R798 vss.n837 vss.n829 251.859
R799 vss.n844 vss 251.859
R800 vss.n832 vss 251.859
R801 vss.n832 vss 251.859
R802 vss.n850 vss.n827 251.859
R803 vss.n839 vss.n827 251.859
R804 vss.n839 vss.n838 251.859
R805 vss.n838 vss.n837 251.859
R806 vss vss.n828 251.859
R807 vss.n845 vss 251.859
R808 vss.n845 vss 251.859
R809 vss vss.n844 251.859
R810 vss.n852 vss.n851 251.859
R811 vss.n851 vss.n850 251.859
R812 vss.n860 vss 251.859
R813 vss vss.n859 251.859
R814 vss.n859 vss 251.859
R815 vss.n828 vss 251.859
R816 vss.n872 vss.n866 251.859
R817 vss.n866 vss.n865 251.859
R818 vss.n865 vss.n822 251.859
R819 vss.n854 vss.n822 251.859
R820 vss vss.n821 251.859
R821 vss vss.n876 251.859
R822 vss.n876 vss 251.859
R823 vss.n860 vss 251.859
R824 vss.n871 vss.n870 251.859
R825 vss.n872 vss.n871 251.859
R826 vss vss.n809 251.859
R827 vss vss.n809 251.859
R828 vss.n821 vss 251.859
R829 vss.n884 vss.n883 251.859
R830 vss.n623 vss.n622 249.667
R831 vss.n929 vss.n203 216.847
R832 vss.n170 vss.n169 213.419
R833 vss.n53 vss.n52 213.407
R834 vss.n887 vss.n886 211.397
R835 vss.n296 vss.n286 209.695
R836 vss.n261 vss.n257 209.695
R837 vss.n972 vss.n971 209.695
R838 vss.n175 vss.n174 209.695
R839 vss.n974 vss.n25 209.695
R840 vss.n110 vss.n39 209.695
R841 vss.n180 vss.n179 209.695
R842 vss.n144 vss.n140 209.695
R843 vss.n372 vss.n339 209.695
R844 vss.n382 vss.n358 209.695
R845 vss.n305 vss.n264 209.695
R846 vss.n331 vss.n330 209.695
R847 vss.n792 vss.n791 188.065
R848 vss.n730 vss.n207 188.065
R849 vss vss.n203 183.087
R850 vss.n932 vss.n931 151.014
R851 vss.n707 vss.n654 150.417
R852 vss.n627 vss.n469 150.417
R853 vss.n523 vss.n518 150.417
R854 vss.n608 vss.n607 150.417
R855 vss.n778 vss.n215 149.835
R856 vss.n778 vss 149.835
R857 vss.n789 vss.n215 149.835
R858 vss.n439 vss.n437 149.835
R859 vss.n439 vss 149.835
R860 vss.n447 vss.n437 149.835
R861 vss.n761 vss.n231 149.835
R862 vss.n761 vss 149.835
R863 vss.n232 vss.n231 149.835
R864 vss.n739 vss.n722 149.835
R865 vss.n739 vss 149.835
R866 vss.n723 vss.n722 149.835
R867 vss.n710 vss.n645 149.835
R868 vss.n710 vss 149.835
R869 vss.n744 vss.n645 149.835
R870 vss.n699 vss.n666 149.835
R871 vss.n679 vss.n671 149.835
R872 vss.n679 vss 149.835
R873 vss.n691 vss.n671 149.835
R874 vss.n675 vss.n672 149.835
R875 vss.n675 vss 149.835
R876 vss.n684 vss.n672 149.835
R877 vss.n732 vss.n726 149.835
R878 vss.n726 vss.n725 149.835
R879 vss.n725 vss 149.835
R880 vss.n716 vss.n715 149.835
R881 vss.n715 vss.n714 149.835
R882 vss.n714 vss 149.835
R883 vss.n502 vss.n487 149.835
R884 vss.n502 vss 149.835
R885 vss.n488 vss.n487 149.835
R886 vss.n512 vss.n477 149.835
R887 vss.n512 vss 149.835
R888 vss.n478 vss.n477 149.835
R889 vss.n615 vss.n614 149.835
R890 vss.n577 vss.n549 149.835
R891 vss.n577 vss 149.835
R892 vss.n594 vss.n549 149.835
R893 vss.n563 vss.n559 149.835
R894 vss.n563 vss 149.835
R895 vss.n574 vss.n559 149.835
R896 vss.n497 vss.n491 149.835
R897 vss.n491 vss.n490 149.835
R898 vss.n490 vss 149.835
R899 vss.n508 vss.n480 149.835
R900 vss.n480 vss.n479 149.835
R901 vss.n479 vss 149.835
R902 vss.n583 vss.n582 149.835
R903 vss.n582 vss.n581 149.835
R904 vss.n581 vss 149.835
R905 vss.n569 vss.n568 149.835
R906 vss.n568 vss.n560 149.835
R907 vss.n560 vss 149.835
R908 vss.n619 vss.n527 149.835
R909 vss.n589 vss.n588 149.835
R910 vss.n765 vss.n222 149.835
R911 vss.n765 vss 149.835
R912 vss.n775 vss.n222 149.835
R913 vss.n784 vss.n783 149.835
R914 vss.n783 vss.n216 149.835
R915 vss.n216 vss 149.835
R916 vss.n225 vss 149.835
R917 vss.n770 vss.n225 149.835
R918 vss.n771 vss.n770 149.835
R919 vss.n789 vss.n788 149.459
R920 vss.n448 vss.n447 149.459
R921 vss.n760 vss.n232 149.459
R922 vss.n738 vss.n723 149.459
R923 vss.n745 vss.n744 149.459
R924 vss.n691 vss.n690 149.459
R925 vss.n685 vss.n684 149.459
R926 vss.n733 vss.n732 149.459
R927 vss.n716 vss.n643 149.459
R928 vss.n501 vss.n488 149.459
R929 vss.n511 vss.n478 149.459
R930 vss.n595 vss.n594 149.459
R931 vss.n574 vss.n573 149.459
R932 vss.n498 vss.n497 149.459
R933 vss.n509 vss.n508 149.459
R934 vss.n583 vss.n548 149.459
R935 vss.n570 vss.n569 149.459
R936 vss.n775 vss.n774 149.459
R937 vss.n785 vss.n784 149.459
R938 vss.n772 vss.n771 149.459
R939 vss.n622 vss.n621 132.8
R940 vss.n608 vss 132.129
R941 vss.n707 vss 132.127
R942 vss vss.n469 132.127
R943 vss vss.n666 130.802
R944 vss.n615 vss 130.802
R945 vss.n589 vss 130.802
R946 vss.n763 vss.n228 125.897
R947 vss.n442 vss.n228 125.897
R948 vss.n444 vss.n443 125.897
R949 vss.n444 vss.n209 125.897
R950 vss.n621 vss.n620 120.001
R951 vss vss 118.966
R952 vss.n935 vss.n202 117.272
R953 vss.n928 vss.n890 117.001
R954 vss.n895 vss.n890 117.001
R955 vss.n896 vss.n891 117.001
R956 vss.n923 vss.n896 117.001
R957 vss.n917 vss 117.001
R958 vss.n917 vss.n916 117.001
R959 vss.n910 vss.n909 117.001
R960 vss.n909 vss.n908 117.001
R961 vss vss.n903 117.001
R962 vss.n915 vss.n899 117.001
R963 vss.n916 vss.n915 117.001
R964 vss.n922 vss 117.001
R965 vss.n923 vss.n922 117.001
R966 vss vss.n889 117.001
R967 vss.n895 vss.n889 117.001
R968 vss.n205 vss.n202 117.001
R969 vss.n204 vss 117.001
R970 vss.n205 vss.n204 117.001
R971 vss.n374 vss.n373 117.001
R972 vss.n375 vss.n374 117.001
R973 vss.n369 vss.n368 117.001
R974 vss.n375 vss.n369 117.001
R975 vss.n400 vss.n399 117.001
R976 vss.n402 vss.n400 117.001
R977 vss.n404 vss.n403 117.001
R978 vss.n403 vss.n402 117.001
R979 vss.n299 vss.n298 117.001
R980 vss.n298 vss.n267 117.001
R981 vss.n240 vss.n238 117.001
R982 vss.n245 vss.n240 117.001
R983 vss.n416 vss.n415 117.001
R984 vss.n415 vss.n245 117.001
R985 vss.n288 vss.n287 117.001
R986 vss.n288 vss.n241 117.001
R987 vss.n292 vss.n291 117.001
R988 vss.n291 vss.n241 117.001
R989 vss.n260 vss.n259 117.001
R990 vss.n411 vss.n259 117.001
R991 vss.n282 vss.n280 117.001
R992 vss.n280 vss.n210 117.001
R993 vss.n285 vss.n284 117.001
R994 vss.n284 vss.n267 117.001
R995 vss.n408 vss.n407 117.001
R996 vss.n409 vss.n408 117.001
R997 vss.n318 vss.n317 117.001
R998 vss.n317 vss.n241 117.001
R999 vss.n315 vss.n263 117.001
R1000 vss.n315 vss.n241 117.001
R1001 vss.n410 vss.n251 117.001
R1002 vss.n411 vss.n410 117.001
R1003 vss.n277 vss.n274 117.001
R1004 vss.n277 vss.n267 117.001
R1005 vss.n273 vss.n272 117.001
R1006 vss.n272 vss.n267 117.001
R1007 vss.n276 vss.n275 117.001
R1008 vss.n276 vss.n210 117.001
R1009 vss.n329 vss.n328 117.001
R1010 vss.n328 vss.n245 117.001
R1011 vss.n424 vss.n248 117.001
R1012 vss.n248 vss.n245 117.001
R1013 vss.n771 vss.n219 117.001
R1014 vss.n777 vss.n219 117.001
R1015 vss.n768 vss.n225 117.001
R1016 vss.n768 vss.n767 117.001
R1017 vss.n784 vss.n212 117.001
R1018 vss.n791 vss.n212 117.001
R1019 vss.n781 vss.n216 117.001
R1020 vss.n781 vss.n780 117.001
R1021 vss.n776 vss.n775 117.001
R1022 vss.n777 vss.n776 117.001
R1023 vss.n766 vss.n765 117.001
R1024 vss.n767 vss.n766 117.001
R1025 vss.n790 vss.n789 117.001
R1026 vss.n791 vss.n790 117.001
R1027 vss.n779 vss.n778 117.001
R1028 vss.n780 vss.n779 117.001
R1029 vss.n441 vss.n232 117.001
R1030 vss.n442 vss.n441 117.001
R1031 vss.n762 vss.n761 117.001
R1032 vss.n763 vss.n762 117.001
R1033 vss.n447 vss.n446 117.001
R1034 vss.n446 vss.n209 117.001
R1035 vss.n440 vss.n439 117.001
R1036 vss.n443 vss.n440 117.001
R1037 vss.n717 vss.n716 117.001
R1038 vss.n742 vss.n717 117.001
R1039 vss.n714 vss.n713 117.001
R1040 vss.n713 vss.n712 117.001
R1041 vss.n732 vss.n731 117.001
R1042 vss.n731 vss.n730 117.001
R1043 vss.n725 vss.n718 117.001
R1044 vss.n741 vss.n718 117.001
R1045 vss.n684 vss.n683 117.001
R1046 vss.n683 vss.n682 117.001
R1047 vss.n676 vss.n675 117.001
R1048 vss.n677 vss.n676 117.001
R1049 vss.n692 vss.n691 117.001
R1050 vss.n693 vss.n692 117.001
R1051 vss.n680 vss.n679 117.001
R1052 vss.n681 vss.n680 117.001
R1053 vss.n665 vss.n664 117.001
R1054 vss.n664 vss.n659 117.001
R1055 vss.n662 vss.n655 117.001
R1056 vss.n662 vss.n660 117.001
R1057 vss.n708 vss.n707 117.001
R1058 vss.n709 vss.n708 117.001
R1059 vss.n667 vss.n666 117.001
R1060 vss.n694 vss.n667 117.001
R1061 vss.n744 vss.n743 117.001
R1062 vss.n743 vss.n742 117.001
R1063 vss.n711 vss.n710 117.001
R1064 vss.n712 vss.n711 117.001
R1065 vss.n729 vss.n723 117.001
R1066 vss.n730 vss.n729 117.001
R1067 vss.n740 vss.n739 117.001
R1068 vss.n741 vss.n740 117.001
R1069 vss.n569 vss.n556 117.001
R1070 vss.n576 vss.n556 117.001
R1071 vss.n566 vss.n560 117.001
R1072 vss.n566 vss.n565 117.001
R1073 vss.n584 vss.n583 117.001
R1074 vss.n592 vss.n584 117.001
R1075 vss.n581 vss.n580 117.001
R1076 vss.n580 vss.n579 117.001
R1077 vss.n546 vss.n545 117.001
R1078 vss.n545 vss.n540 117.001
R1079 vss.n543 vss.n536 117.001
R1080 vss.n543 vss.n541 117.001
R1081 vss.n609 vss.n608 117.001
R1082 vss.n610 vss.n609 117.001
R1083 vss.n590 vss.n589 117.001
R1084 vss.n591 vss.n590 117.001
R1085 vss.n530 vss.n522 117.001
R1086 vss.n530 vss.n458 117.001
R1087 vss.n521 vss.n520 117.001
R1088 vss.n520 vss.n460 117.001
R1089 vss.n518 vss.n517 117.001
R1090 vss.n517 vss.n515 117.001
R1091 vss.n619 vss.n618 117.001
R1092 vss.n618 vss.n617 117.001
R1093 vss.n508 vss.n507 117.001
R1094 vss.n507 vss.n506 117.001
R1095 vss.n479 vss.n473 117.001
R1096 vss.n514 vss.n473 117.001
R1097 vss.n497 vss.n496 117.001
R1098 vss.n496 vss.n495 117.001
R1099 vss.n490 vss.n483 117.001
R1100 vss.n504 vss.n483 117.001
R1101 vss.n575 vss.n574 117.001
R1102 vss.n576 vss.n575 117.001
R1103 vss.n564 vss.n563 117.001
R1104 vss.n565 vss.n564 117.001
R1105 vss.n594 vss.n593 117.001
R1106 vss.n593 vss.n592 117.001
R1107 vss.n578 vss.n577 117.001
R1108 vss.n579 vss.n578 117.001
R1109 vss.n465 vss.n464 117.001
R1110 vss.n464 vss.n458 117.001
R1111 vss.n468 vss.n467 117.001
R1112 vss.n467 vss.n460 117.001
R1113 vss.n470 vss.n469 117.001
R1114 vss.n515 vss.n470 117.001
R1115 vss.n616 vss.n615 117.001
R1116 vss.n617 vss.n616 117.001
R1117 vss.n505 vss.n478 117.001
R1118 vss.n506 vss.n505 117.001
R1119 vss.n513 vss.n512 117.001
R1120 vss.n514 vss.n513 117.001
R1121 vss.n494 vss.n488 117.001
R1122 vss.n495 vss.n494 117.001
R1123 vss.n503 vss.n502 117.001
R1124 vss.n504 vss.n503 117.001
R1125 vss.n383 vss.n361 117.001
R1126 vss.n388 vss.n361 117.001
R1127 vss.n390 vss.n389 117.001
R1128 vss.n389 vss.n388 117.001
R1129 vss.n365 vss.n364 117.001
R1130 vss.n365 vss.n362 117.001
R1131 vss.n984 vss.n983 117.001
R1132 vss.n983 vss.n982 117.001
R1133 vss.n105 vss.n66 117.001
R1134 vss.n964 vss.n66 117.001
R1135 vss.n107 vss.n28 117.001
R1136 vss.n982 vss.n28 117.001
R1137 vss.n959 vss.n62 117.001
R1138 vss.n964 vss.n62 117.001
R1139 vss.n981 vss.n980 117.001
R1140 vss.n982 vss.n981 117.001
R1141 vss.n111 vss.n34 117.001
R1142 vss.n982 vss.n34 117.001
R1143 vss.n22 vss.n20 117.001
R1144 vss.n982 vss.n20 117.001
R1145 vss.n963 vss.n23 117.001
R1146 vss.n964 vss.n963 117.001
R1147 vss.n970 vss.n33 117.001
R1148 vss.n982 vss.n33 117.001
R1149 vss.n120 vss.n63 117.001
R1150 vss.n964 vss.n63 117.001
R1151 vss.n114 vss.n64 117.001
R1152 vss.n964 vss.n64 117.001
R1153 vss.n50 vss.n30 117.001
R1154 vss.n982 vss.n30 117.001
R1155 vss.n51 vss.n32 117.001
R1156 vss.n982 vss.n32 117.001
R1157 vss.n49 vss.n29 117.001
R1158 vss.n982 vss.n29 117.001
R1159 vss.n966 vss.n965 117.001
R1160 vss.n965 vss.n964 117.001
R1161 vss.n178 vss.n131 117.001
R1162 vss.n188 vss.n131 117.001
R1163 vss.n139 vss.n132 117.001
R1164 vss.n188 vss.n132 117.001
R1165 vss.n143 vss.n136 117.001
R1166 vss.n188 vss.n136 117.001
R1167 vss.n187 vss.n186 117.001
R1168 vss.n188 vss.n187 117.001
R1169 vss.n93 vss.n92 117.001
R1170 vss.n92 vss.n76 117.001
R1171 vss.n75 vss.n73 117.001
R1172 vss.n76 vss.n75 117.001
R1173 vss.n950 vss.n79 117.001
R1174 vss.n79 vss.n76 117.001
R1175 vss.n82 vss.n81 117.001
R1176 vss.n188 vss.n82 117.001
R1177 vss.n152 vss.n135 117.001
R1178 vss.n188 vss.n135 117.001
R1179 vss.n189 vss.n129 117.001
R1180 vss.n189 vss.n188 117.001
R1181 vss.n168 vss.n134 117.001
R1182 vss.n188 vss.n134 117.001
R1183 vss.n156 vss.n155 117.001
R1184 vss.n155 vss.n76 117.001
R1185 vss.n192 vss.n191 117.001
R1186 vss.n191 vss.n76 117.001
R1187 vss.n160 vss.n159 117.001
R1188 vss.n159 vss.n76 117.001
R1189 vss.n151 vss.n133 117.001
R1190 vss.n188 vss.n133 117.001
R1191 vss vss.n452 115.576
R1192 vss.n907 vss.n903 109.642
R1193 vss.n793 vss.n210 108.163
R1194 vss.n946 vss.n76 101.77
R1195 vss.n953 vss.n76 101.77
R1196 vss.n964 vss.n61 101.77
R1197 vss.n964 vss.n13 100.514
R1198 vss.n931 vss.n888 96.1003
R1199 vss.n401 vss.n336 90.9521
R1200 vss.n701 vss.n655 90.3534
R1201 vss.n706 vss.n655 90.3534
R1202 vss.n700 vss.n665 90.3534
R1203 vss.n695 vss.n665 90.3534
R1204 vss.n628 vss.n468 90.3534
R1205 vss.n468 vss.n455 90.3534
R1206 vss.n466 vss.n465 90.3534
R1207 vss.n465 vss.n454 90.3534
R1208 vss.n620 vss.n522 90.3534
R1209 vss.n526 vss.n522 90.3534
R1210 vss.n622 vss.n521 90.3534
R1211 vss.n524 vss.n521 90.3534
R1212 vss.n547 vss.n546 90.3534
R1213 vss.n546 vss.n537 90.3534
R1214 vss.n601 vss.n536 90.3534
R1215 vss.n606 vss.n536 90.3534
R1216 vss.n623 vss.n518 89.9911
R1217 vss.n976 vss.n31 89.6255
R1218 vss vss.n904 89.224
R1219 vss vss.n900 89.224
R1220 vss.n911 vss 89.224
R1221 vss.n911 vss.n910 89.224
R1222 vss vss.n892 89.224
R1223 vss vss.n921 89.224
R1224 vss.n921 vss.n899 89.224
R1225 vss.n904 vss.n899 89.224
R1226 vss.n892 vss 89.224
R1227 vss.n928 vss.n927 89.224
R1228 vss.n927 vss.n891 89.224
R1229 vss.n900 vss.n891 89.224
R1230 vss.n87 vss.n4 86.561
R1231 vss.n182 vss.n130 86.275
R1232 vss.n287 vss.n237 85.0829
R1233 vss.n287 vss.n255 85.0829
R1234 vss.n294 vss.n292 85.0829
R1235 vss.n416 vss.n257 85.0829
R1236 vss.n299 vss.n296 85.0829
R1237 vss.n55 vss.n50 85.0829
R1238 vss.n53 vss.n51 85.0829
R1239 vss.n971 vss.n970 85.0829
R1240 vss.n115 vss.n114 85.0829
R1241 vss.n114 vss.n9 85.0829
R1242 vss.n172 vss.n168 85.0829
R1243 vss.n167 vss.n156 85.0829
R1244 vss.n156 vss.n126 85.0829
R1245 vss.n174 vss.n152 85.0829
R1246 vss.n170 vss.n129 85.0829
R1247 vss.n107 vss.n39 85.0829
R1248 vss.n984 vss.n25 85.0829
R1249 vss.n960 vss.n959 85.0829
R1250 vss.n959 vss.n37 85.0829
R1251 vss.n980 vss.n979 85.0829
R1252 vss.n186 vss.n185 85.0829
R1253 vss.n94 vss.n93 85.0829
R1254 vss.n93 vss.n72 85.0829
R1255 vss.n179 vss.n178 85.0829
R1256 vss.n140 vss.n139 85.0829
R1257 vss.n368 vss.n367 85.0829
R1258 vss.n399 vss.n347 85.0829
R1259 vss.n399 vss.n398 85.0829
R1260 vss.n373 vss.n372 85.0829
R1261 vss.n383 vss.n382 85.0829
R1262 vss.n318 vss.n314 85.0829
R1263 vss.n319 vss.n318 85.0829
R1264 vss.n325 vss.n263 85.0829
R1265 vss.n274 vss.n264 85.0829
R1266 vss.n330 vss.n329 85.0829
R1267 vss.n303 vss.n282 84.9588
R1268 vss.n57 vss.n49 84.9588
R1269 vss.n161 vss.n151 84.9588
R1270 vss.n987 vss.n22 84.9588
R1271 vss.n948 vss.n81 84.9588
R1272 vss.n407 vss.n406 84.9588
R1273 vss.n309 vss.n275 84.9588
R1274 vss.n422 vss.n251 84.6953
R1275 vss.n260 vss.n252 84.6953
R1276 vss.n143 vss.n104 84.6953
R1277 vss.n112 vss.n111 84.6953
R1278 vss.n391 vss.n390 84.6953
R1279 vss.n946 vss.n87 83.5719
R1280 vss.n443 vss.n442 82.869
R1281 vss vss.n623 77.2563
R1282 vss.n982 vss.n27 71.1979
R1283 vss.n300 vss.n255 66.6518
R1284 vss.n968 vss.n9 66.6518
R1285 vss.n167 vss.n164 66.6518
R1286 vss.n37 vss.n24 66.6518
R1287 vss.n96 vss.n94 66.6518
R1288 vss.n353 vss.n347 66.6518
R1289 vss.n314 vss.n312 66.6518
R1290 vss.n418 vss.n417 64.7759
R1291 vss.n166 vss.n165 64.7759
R1292 vss.n991 vss.n10 64.7759
R1293 vss.n108 vss.n106 64.7759
R1294 vss.n944 vss.n95 64.7759
R1295 vss.n385 vss.n384 64.7759
R1296 vss.n313 vss.n249 64.7759
R1297 vss.n188 vss.n27 64.497
R1298 vss.n418 vss.n255 63.1207
R1299 vss.n167 vss.n166 63.1207
R1300 vss.n991 vss.n9 63.1207
R1301 vss.n106 vss.n37 63.1207
R1302 vss.n944 vss.n94 63.1207
R1303 vss.n385 vss.n347 63.1207
R1304 vss.n314 vss.n313 63.1207
R1305 vss.n301 vss.n300 61.2449
R1306 vss.n969 vss.n968 61.2449
R1307 vss.n164 vss.n163 61.2449
R1308 vss.n985 vss.n24 61.2449
R1309 vss.n96 vss.n80 61.2449
R1310 vss.n353 vss.n340 61.2449
R1311 vss.n312 vss.n311 61.2449
R1312 vss.n700 vss.n699 59.4829
R1313 vss.n702 vss.n700 59.4829
R1314 vss.n702 vss.n701 59.4829
R1315 vss.n701 vss.n654 59.4829
R1316 vss.n614 vss.n466 59.4829
R1317 vss.n629 vss.n466 59.4829
R1318 vss.n629 vss.n628 59.4829
R1319 vss.n628 vss.n627 59.4829
R1320 vss.n527 vss.n526 59.4829
R1321 vss.n526 vss.n525 59.4829
R1322 vss.n525 vss.n524 59.4829
R1323 vss.n524 vss.n523 59.4829
R1324 vss.n588 vss.n537 59.4829
R1325 vss.n605 vss.n537 59.4829
R1326 vss.n606 vss.n605 59.4829
R1327 vss.n607 vss.n606 59.4829
R1328 vss.n417 vss.n416 58.5793
R1329 vss.n301 vss.n299 58.5793
R1330 vss.n51 vss.n10 58.5793
R1331 vss.n970 vss.n969 58.5793
R1332 vss.n163 vss.n152 58.5793
R1333 vss.n165 vss.n129 58.5793
R1334 vss.n108 vss.n107 58.5793
R1335 vss.n985 vss.n984 58.5793
R1336 vss.n178 vss.n80 58.5793
R1337 vss.n139 vss.n95 58.5793
R1338 vss.n373 vss.n340 58.5793
R1339 vss.n384 vss.n383 58.5793
R1340 vss.n311 vss.n274 58.5793
R1341 vss.n329 vss.n249 58.5793
R1342 vss.n292 vss.n255 54.2123
R1343 vss.n50 vss.n9 54.2123
R1344 vss.n168 vss.n167 54.2123
R1345 vss.n980 vss.n37 54.2123
R1346 vss.n186 vss.n94 54.2123
R1347 vss.n368 vss.n347 54.2123
R1348 vss.n314 vss.n263 54.2123
R1349 vss.n794 vss.n209 42.2316
R1350 vss.n406 vss.n338 41.7862
R1351 vss.n344 vss.n338 41.7862
R1352 vss.n339 vss.n337 41.7862
R1353 vss.n376 vss.n337 41.7862
R1354 vss.n333 vss.n252 41.7862
R1355 vss.n412 vss.n333 41.7862
R1356 vss.n413 vss.n261 41.7862
R1357 vss.n413 vss.n412 41.7862
R1358 vss.n286 vss.n279 41.7862
R1359 vss.n307 vss.n279 41.7862
R1360 vss.n304 vss.n303 41.7862
R1361 vss.n307 vss.n304 41.7862
R1362 vss.n309 vss.n308 41.7862
R1363 vss.n308 vss.n307 41.7862
R1364 vss.n306 vss.n305 41.7862
R1365 vss.n307 vss.n306 41.7862
R1366 vss.n332 vss.n331 41.7862
R1367 vss.n412 vss.n332 41.7862
R1368 vss.n422 vss.n250 41.7862
R1369 vss.n412 vss.n250 41.7862
R1370 vss.n391 vss.n357 41.7862
R1371 vss.n387 vss.n357 41.7862
R1372 vss.n359 vss.n358 41.7862
R1373 vss.n360 vss.n359 41.7862
R1374 vss.n112 vss.n15 41.7862
R1375 vss.n989 vss.n15 41.7862
R1376 vss.n110 vss.n42 41.7862
R1377 vss.n976 vss.n42 41.7862
R1378 vss.n975 vss.n974 41.7862
R1379 vss.n976 vss.n975 41.7862
R1380 vss.n988 vss.n987 41.7862
R1381 vss.n989 vss.n988 41.7862
R1382 vss.n976 vss.n44 41.7862
R1383 vss.n973 vss.n972 41.7862
R1384 vss.n976 vss.n973 41.7862
R1385 vss.n57 vss.n18 41.7862
R1386 vss.n989 vss.n18 41.7862
R1387 vss.n104 vss.n85 41.7862
R1388 vss.n946 vss.n85 41.7862
R1389 vss.n948 vss.n947 41.7862
R1390 vss.n947 vss.n946 41.7862
R1391 vss.n181 vss.n180 41.7862
R1392 vss.n182 vss.n181 41.7862
R1393 vss.n145 vss.n144 41.7862
R1394 vss.n182 vss.n145 41.7862
R1395 vss.n161 vss.n89 41.7862
R1396 vss.n946 vss.n89 41.7862
R1397 vss.n176 vss.n175 41.7862
R1398 vss.n182 vss.n176 41.7862
R1399 vss.n182 vss.n147 41.7862
R1400 vss.n127 vss.n4 41.0949
R1401 vss vss.n695 40.4485
R1402 vss.n706 vss 40.4485
R1403 vss vss.n706 40.4485
R1404 vss vss.n454 40.4485
R1405 vss vss.n455 40.4485
R1406 vss vss.n455 40.4485
R1407 vss vss.n547 40.4485
R1408 vss vss.n601 40.4485
R1409 vss.n601 vss 40.4485
R1410 vss.n695 vss.n656 38.1445
R1411 vss.n633 vss.n454 38.1445
R1412 vss.n600 vss.n547 38.1445
R1413 vss.n52 vss.n44 37.7132
R1414 vss.n169 vss.n147 37.6975
R1415 vss.n946 vss.n27 37.2744
R1416 vss.n934 vss.n933 34.4123
R1417 vss.n933 vss.n932 34.4123
R1418 vss.n334 vss.n201 34.4123
R1419 vss.n335 vss.n334 34.4123
R1420 vss.n353 vss.n352 34.4123
R1421 vss.n352 vss.n344 34.4123
R1422 vss.n343 vss.n341 34.4123
R1423 vss.n401 vss.n343 34.4123
R1424 vss.n377 vss.n371 34.4123
R1425 vss.n377 vss.n376 34.4123
R1426 vss.n300 vss.n270 34.4123
R1427 vss.n322 vss.n270 34.4123
R1428 vss.n418 vss.n244 34.4123
R1429 vss.n427 vss.n244 34.4123
R1430 vss.n293 vss.n246 34.4123
R1431 vss.n427 vss.n246 34.4123
R1432 vss.n295 vss.n271 34.4123
R1433 vss.n322 vss.n271 34.4123
R1434 vss.n283 vss.n269 34.4123
R1435 vss.n322 vss.n269 34.4123
R1436 vss.n429 vss.n428 34.4123
R1437 vss.n428 vss.n427 34.4123
R1438 vss.n426 vss.n425 34.4123
R1439 vss.n427 vss.n426 34.4123
R1440 vss.n321 vss.n320 34.4123
R1441 vss.n322 vss.n321 34.4123
R1442 vss.n312 vss.n268 34.4123
R1443 vss.n322 vss.n268 34.4123
R1444 vss.n313 vss.n243 34.4123
R1445 vss.n427 vss.n243 34.4123
R1446 vss.n324 vss.n323 34.4123
R1447 vss.n323 vss.n322 34.4123
R1448 vss.n326 vss.n242 34.4123
R1449 vss.n427 vss.n242 34.4123
R1450 vss.n386 vss.n385 34.4123
R1451 vss.n387 vss.n386 34.4123
R1452 vss.n363 vss.n348 34.4123
R1453 vss.n363 vss.n206 34.4123
R1454 vss.n381 vss.n380 34.4123
R1455 vss.n380 vss.n360 34.4123
R1456 vss.n24 vss.n14 34.4123
R1457 vss.n989 vss.n14 34.4123
R1458 vss.n106 vss.n19 34.4123
R1459 vss.n989 vss.n19 34.4123
R1460 vss.n978 vss.n977 34.4123
R1461 vss.n977 vss.n976 34.4123
R1462 vss.n41 vss.n38 34.4123
R1463 vss.n976 vss.n41 34.4123
R1464 vss.n962 vss.n961 34.4123
R1465 vss.n962 vss.n61 34.4123
R1466 vss.n69 vss.n68 34.4123
R1467 vss.n68 vss.n61 34.4123
R1468 vss.n968 vss.n16 34.4123
R1469 vss.n989 vss.n16 34.4123
R1470 vss.n991 vss.n990 34.4123
R1471 vss.n990 vss.n989 34.4123
R1472 vss.n54 vss.n47 34.4123
R1473 vss.n976 vss.n47 34.4123
R1474 vss.n56 vss.n43 34.4123
R1475 vss.n976 vss.n43 34.4123
R1476 vss.n59 vss.n58 34.4123
R1477 vss.n61 vss.n59 34.4123
R1478 vss.n123 vss.n122 34.4123
R1479 vss.n122 vss.n61 34.4123
R1480 vss.n96 vss.n84 34.4123
R1481 vss.n946 vss.n84 34.4123
R1482 vss.n945 vss.n944 34.4123
R1483 vss.n946 vss.n945 34.4123
R1484 vss.n955 vss.n954 34.4123
R1485 vss.n954 vss.n953 34.4123
R1486 vss.n952 vss.n951 34.4123
R1487 vss.n953 vss.n952 34.4123
R1488 vss.n142 vss.n138 34.4123
R1489 vss.n182 vss.n142 34.4123
R1490 vss.n184 vss.n183 34.4123
R1491 vss.n183 vss.n182 34.4123
R1492 vss.n164 vss.n86 34.4123
R1493 vss.n946 vss.n86 34.4123
R1494 vss.n166 vss.n88 34.4123
R1495 vss.n946 vss.n88 34.4123
R1496 vss.n193 vss.n77 34.4123
R1497 vss.n953 vss.n77 34.4123
R1498 vss.n157 vss.n78 34.4123
R1499 vss.n953 vss.n78 34.4123
R1500 vss.n173 vss.n146 34.4123
R1501 vss.n182 vss.n146 34.4123
R1502 vss.n171 vss.n149 34.4123
R1503 vss.n182 vss.n149 34.4123
R1504 vss.n829 vss.n799 32.5005
R1505 vss.n886 vss.n799 32.5005
R1506 vss vss.n816 32.5005
R1507 vss.n878 vss.n816 32.5005
R1508 vss vss.n815 32.5005
R1509 vss.n878 vss.n815 32.5005
R1510 vss.n838 vss.n801 32.5005
R1511 vss.n886 vss.n801 32.5005
R1512 vss vss.n814 32.5005
R1513 vss.n878 vss.n814 32.5005
R1514 vss.n851 vss.n802 32.5005
R1515 vss.n886 vss.n802 32.5005
R1516 vss.n827 vss.n798 32.5005
R1517 vss.n886 vss.n798 32.5005
R1518 vss vss.n817 32.5005
R1519 vss.n878 vss.n817 32.5005
R1520 vss.n853 vss.n797 32.5005
R1521 vss.n886 vss.n797 32.5005
R1522 vss vss.n818 32.5005
R1523 vss.n878 vss.n818 32.5005
R1524 vss vss.n813 32.5005
R1525 vss.n878 vss.n813 32.5005
R1526 vss.n822 vss.n803 32.5005
R1527 vss.n886 vss.n803 32.5005
R1528 vss vss.n812 32.5005
R1529 vss.n878 vss.n812 32.5005
R1530 vss.n871 vss.n804 32.5005
R1531 vss.n886 vss.n804 32.5005
R1532 vss.n866 vss.n796 32.5005
R1533 vss.n886 vss.n796 32.5005
R1534 vss.n877 vss 32.5005
R1535 vss.n878 vss.n877 32.5005
R1536 vss.n808 vss.n795 32.5005
R1537 vss.n886 vss.n795 32.5005
R1538 vss.n879 vss 32.5005
R1539 vss.n879 vss.n878 32.5005
R1540 vss vss.n810 32.5005
R1541 vss.n878 vss.n810 32.5005
R1542 vss.n885 vss.n884 32.5005
R1543 vss.n886 vss.n885 32.5005
R1544 vss.n27 vss.n17 24.7102
R1545 vss.n887 vss.n61 22.1973
R1546 vss.n831 vss.n830 19.5005
R1547 vss.n830 vss.n800 19.5005
R1548 vss.n836 vss.n835 19.5005
R1549 vss.n835 vss.n800 19.5005
R1550 vss.n843 vss.n842 19.5005
R1551 vss.n842 vss.n800 19.5005
R1552 vss.n849 vss.n848 19.5005
R1553 vss.n848 vss.n800 19.5005
R1554 vss.n826 vss.n825 19.5005
R1555 vss.n825 vss.n800 19.5005
R1556 vss.n858 vss.n857 19.5005
R1557 vss.n857 vss.n800 19.5005
R1558 vss.n864 vss.n863 19.5005
R1559 vss.n863 vss.n800 19.5005
R1560 vss.n875 vss.n874 19.5005
R1561 vss.n874 vss.n800 19.5005
R1562 vss.n869 vss.n868 19.5005
R1563 vss.n868 vss.n800 19.5005
R1564 vss.n882 vss.n881 19.5005
R1565 vss.n881 vss.n800 19.5005
R1566 vss.n807 vss.n805 19.5005
R1567 vss.n805 vss.n800 19.5005
R1568 vss.n953 vss.n27 18.8469
R1569 vss.n417 vss.n256 18.297
R1570 vss.n302 vss.n301 18.297
R1571 vss.n119 vss.n10 18.297
R1572 vss.n969 vss.n967 18.297
R1573 vss.n163 vss.n162 18.297
R1574 vss.n165 vss.n127 18.297
R1575 vss.n109 vss.n108 18.297
R1576 vss.n986 vss.n985 18.297
R1577 vss.n949 vss.n80 18.297
R1578 vss.n103 vss.n95 18.297
R1579 vss.n405 vss.n340 18.297
R1580 vss.n384 vss.n356 18.297
R1581 vss.n311 vss.n310 18.297
R1582 vss.n423 vss.n249 18.297
R1583 vss.n926 vss.n925 17.2064
R1584 vss.n925 vss.n924 17.2064
R1585 vss.n920 vss.n919 17.2064
R1586 vss.n919 vss.n897 17.2064
R1587 vss.n913 vss.n912 17.2064
R1588 vss.n913 vss.n902 17.2064
R1589 vss.n906 vss.n905 17.2064
R1590 vss.n930 vss.n929 17.2064
R1591 vss.n931 vss.n930 17.2064
R1592 vss.n188 vss.n130 15.4964
R1593 vss.n994 vss.n4 15.4704
R1594 vss.n982 vss.n31 12.1459
R1595 vss.n303 vss.n302 8.08353
R1596 vss.n256 vss.n252 8.08353
R1597 vss.n967 vss.n57 8.08353
R1598 vss.n162 vss.n161 8.08353
R1599 vss.n987 vss.n986 8.08353
R1600 vss.n112 vss.n109 8.08353
R1601 vss.n949 vss.n948 8.08353
R1602 vss.n104 vss.n103 8.08353
R1603 vss.n406 vss.n405 8.08353
R1604 vss.n391 vss.n356 8.08353
R1605 vss.n310 vss.n309 8.08353
R1606 vss.n423 vss.n422 8.08353
R1607 vss.n758 vss.n757 6.69613
R1608 vss.n989 vss.n17 5.86382
R1609 vss.n908 vss.n907 5.84938
R1610 vss.n636 vss.n451 5.57706
R1611 vss.n642 vss 5.02361
R1612 vss.n453 vss 5.02361
R1613 vss.n453 vss 5.02361
R1614 vss.n598 vss 5.02361
R1615 vss.n450 vss 5.01717
R1616 vss.n436 vss 5.01717
R1617 vss.n687 vss 5.01717
R1618 vss.n688 vss 5.01717
R1619 vss.n644 vss 5.01717
R1620 vss.n644 vss 5.01717
R1621 vss.n736 vss 5.01717
R1622 vss.n736 vss 5.01717
R1623 vss.n571 vss 5.01717
R1624 vss.n571 vss 5.01717
R1625 vss.n597 vss 5.01717
R1626 vss.n597 vss 5.01717
R1627 vss.n489 vss 5.01717
R1628 vss.n489 vss 5.01717
R1629 vss.n499 vss 5.01717
R1630 vss.n499 vss 5.01717
R1631 vss.n223 vss 5.01717
R1632 vss.n223 vss 5.01717
R1633 vss.n786 vss 5.01717
R1634 vss.n786 vss 5.01717
R1635 vss.n686 vss.n638 4.99245
R1636 vss.n735 vss.n734 4.87797
R1637 vss.n724 vss.n641 4.50893
R1638 vss.n751 vss.n639 4.5005
R1639 vss.n753 vss.n752 4.5005
R1640 vss.n748 vss.n747 4.5005
R1641 vss.n734 vss 4.5005
R1642 vss vss.n638 4.5005
R1643 vss.n118 vss.n5 4.3205
R1644 vss.n992 vss.n8 3.27485
R1645 vss.n102 vss.n101 3.27485
R1646 vss.n943 vss.n97 3.27485
R1647 vss.n254 vss.n234 3.27485
R1648 vss.n419 vss.n233 3.27485
R1649 vss.n113 vss.n6 3.27485
R1650 vss.n355 vss.n354 3.27485
R1651 vss.n119 vss.n118 3.24353
R1652 vss.n256 vss.n238 3.08756
R1653 vss.n302 vss.n285 3.08756
R1654 vss.n120 vss.n119 3.08756
R1655 vss.n967 vss.n966 3.08756
R1656 vss.n162 vss.n160 3.08756
R1657 vss.n192 vss.n127 3.08756
R1658 vss.n109 vss.n105 3.08756
R1659 vss.n986 vss.n23 3.08756
R1660 vss.n950 vss.n949 3.08756
R1661 vss.n103 vss.n73 3.08756
R1662 vss.n405 vss.n404 3.08756
R1663 vss.n364 vss.n356 3.08756
R1664 vss.n310 vss.n273 3.08756
R1665 vss.n424 vss.n423 3.08756
R1666 vss.n197 vss 3.06629
R1667 vss.n99 vss 3.06629
R1668 vss.n433 vss 3.06629
R1669 vss.n621 vss 3.01226
R1670 vss.n887 vss.n27 2.6242
R1671 vss.n0 vss 2.51601
R1672 vss.n756 vss.n224 2.46929
R1673 vss.n811 vss.n807 2.35839
R1674 vss vss.n656 2.3045
R1675 vss.n633 vss 2.3045
R1676 vss vss.n600 2.3045
R1677 vss.n0 vss 2.11902
R1678 vss.n994 vss.n5 1.92736
R1679 vss.n236 vss 1.91991
R1680 vss.n125 vss 1.91991
R1681 vss.n71 vss 1.91991
R1682 vss.n760 vss.n759 1.8605
R1683 vss.n449 vss.n448 1.8605
R1684 vss.n746 vss.n643 1.8605
R1685 vss.n737 vss.n733 1.8605
R1686 vss.n686 vss.n685 1.8605
R1687 vss.n690 vss.n689 1.8605
R1688 vss.n746 vss.n745 1.8605
R1689 vss.n738 vss.n737 1.8605
R1690 vss.n572 vss.n570 1.8605
R1691 vss.n596 vss.n548 1.8605
R1692 vss.n510 vss.n509 1.8605
R1693 vss.n500 vss.n498 1.8605
R1694 vss.n573 vss.n572 1.8605
R1695 vss.n596 vss.n595 1.8605
R1696 vss.n511 vss.n510 1.8605
R1697 vss.n501 vss.n500 1.8605
R1698 vss.n787 vss.n785 1.8605
R1699 vss.n774 vss.n773 1.8605
R1700 vss.n788 vss.n787 1.8605
R1701 vss.n773 vss.n772 1.8605
R1702 vss.n637 vss.n636 1.79344
R1703 vss.n993 vss.n6 1.55665
R1704 vss.n993 vss.n992 1.55665
R1705 vss.n942 vss.n102 1.55665
R1706 vss.n943 vss.n942 1.55665
R1707 vss.n393 vss.n355 1.55665
R1708 vss.n420 vss.n254 1.55665
R1709 vss.n420 vss.n419 1.55665
R1710 vss.n198 vss.n113 1.43327
R1711 vss.n198 vss.n8 1.43327
R1712 vss.n101 vss.n100 1.43327
R1713 vss.n100 vss.n97 1.43327
R1714 vss.n354 vss.n200 1.43327
R1715 vss.n434 vss.n234 1.43327
R1716 vss.n434 vss.n233 1.43327
R1717 vss.n940 vss.n939 1.26772
R1718 vss.n989 vss.n13 1.25692
R1719 vss.n936 vss.n201 1.21955
R1720 vss.n757 vss.n756 1.06966
R1721 vss.n749 vss.n748 0.99175
R1722 vss.n420 vss 0.946224
R1723 vss.n993 vss 0.946224
R1724 vss.n942 vss 0.946224
R1725 vss.n432 vss 0.905763
R1726 vss.n196 vss 0.905763
R1727 vss.n70 vss 0.905763
R1728 vss.n941 vss.n104 0.846996
R1729 vss.n941 vss.n112 0.846996
R1730 vss.n392 vss.n391 0.846996
R1731 vss.n422 vss.n421 0.846996
R1732 vss.n421 vss.n252 0.846996
R1733 vss vss 0.771099
R1734 vss.n656 vss.n640 0.715885
R1735 vss.n600 vss.n599 0.715885
R1736 vss.n634 vss.n452 0.715885
R1737 vss.n634 vss.n633 0.715885
R1738 vss.n395 vss 0.695143
R1739 vss.n166 vss.n6 0.664786
R1740 vss.n164 vss.n113 0.664786
R1741 vss.n992 vss.n991 0.664786
R1742 vss.n968 vss.n8 0.664786
R1743 vss.n106 vss.n102 0.664786
R1744 vss.n101 vss.n24 0.664786
R1745 vss.n944 vss.n943 0.664786
R1746 vss.n97 vss.n96 0.664786
R1747 vss.n385 vss.n355 0.664786
R1748 vss.n354 vss.n353 0.664786
R1749 vss.n938 vss 0.664786
R1750 vss.n313 vss.n254 0.664786
R1751 vss.n312 vss.n234 0.664786
R1752 vss.n419 vss.n418 0.664786
R1753 vss.n300 vss.n233 0.664786
R1754 vss.n351 vss 0.644695
R1755 vss vss 0.635531
R1756 vss.n934 vss.n203 0.582318
R1757 vss.n755 vss.n754 0.568833
R1758 vss.n996 vss.n3 0.52089
R1759 vss.n937 vss.n936 0.517167
R1760 vss vss 0.457722
R1761 vss.n253 vss 0.447211
R1762 vss.n7 vss 0.447211
R1763 vss.n98 vss 0.447211
R1764 vss.n100 vss 0.439349
R1765 vss.n198 vss 0.439349
R1766 vss.n434 vss 0.439349
R1767 vss.n749 vss.n639 0.418469
R1768 vss.n751 vss.n750 0.418469
R1769 vss.n754 vss.n753 0.414451
R1770 vss vss 0.406319
R1771 vss.n599 vss 0.405187
R1772 vss.n635 vss.n634 0.402844
R1773 vss.n750 vss.n640 0.401281
R1774 vss.n788 vss 0.376971
R1775 vss.n448 vss 0.376971
R1776 vss vss.n760 0.376971
R1777 vss.n430 vss.n237 0.376971
R1778 vss.n124 vss.n115 0.376971
R1779 vss.n194 vss.n126 0.376971
R1780 vss.n960 vss.n958 0.376971
R1781 vss.n956 vss.n72 0.376971
R1782 vss.n398 vss.n397 0.376971
R1783 vss.n319 vss.n235 0.376971
R1784 vss vss.n738 0.376971
R1785 vss.n745 vss 0.376971
R1786 vss.n690 vss 0.376971
R1787 vss.n685 vss 0.376971
R1788 vss.n733 vss 0.376971
R1789 vss vss.n643 0.376971
R1790 vss vss.n501 0.376971
R1791 vss vss.n511 0.376971
R1792 vss.n595 vss 0.376971
R1793 vss.n573 vss 0.376971
R1794 vss.n498 vss 0.376971
R1795 vss.n509 vss 0.376971
R1796 vss vss.n548 0.376971
R1797 vss.n570 vss 0.376971
R1798 vss.n621 vss.n452 0.376971
R1799 vss.n774 vss 0.376971
R1800 vss.n785 vss 0.376971
R1801 vss.n772 vss 0.376971
R1802 vss.n642 vss.n640 0.376281
R1803 vss.n599 vss.n598 0.376281
R1804 vss.n634 vss.n453 0.376281
R1805 vss.n748 vss.n641 0.35393
R1806 vss.n435 vss.n434 0.346566
R1807 vss.n393 vss 0.342762
R1808 vss.n253 vss.n236 0.321553
R1809 vss.n433 vss.n432 0.321553
R1810 vss.n125 vss.n7 0.321553
R1811 vss.n197 vss.n196 0.321553
R1812 vss.n98 vss.n71 0.321553
R1813 vss.n99 vss.n70 0.321553
R1814 vss.n394 vss 0.318384
R1815 vss.n811 vss.n2 0.304262
R1816 vss.n753 vss.n639 0.301281
R1817 vss.n752 vss.n751 0.301281
R1818 vss.n755 vss.n637 0.250766
R1819 vss.n756 vss.n755 0.250595
R1820 vss.n395 vss.n394 0.228964
R1821 vss.n997 vss.n2 0.222309
R1822 vss.n2 vss.n1 0.218382
R1823 vss vss.n449 0.208833
R1824 vss.n1 vss.n0 0.188289
R1825 vss.n432 vss.n431 0.186355
R1826 vss.n196 vss.n195 0.186355
R1827 vss.n957 vss.n70 0.186355
R1828 vss.n996 vss.n995 0.181262
R1829 vss.n420 vss.n253 0.171553
R1830 vss.n993 vss.n7 0.171553
R1831 vss.n942 vss.n98 0.171553
R1832 vss.n199 vss 0.166889
R1833 vss vss.n746 0.166125
R1834 vss.n510 vss 0.166125
R1835 vss.n689 vss 0.164562
R1836 vss.n737 vss 0.164562
R1837 vss.n596 vss 0.164562
R1838 vss.n500 vss 0.164562
R1839 vss.n787 vss 0.164562
R1840 vss.n431 vss.n236 0.158395
R1841 vss.n195 vss.n125 0.158395
R1842 vss.n957 vss.n71 0.158395
R1843 vss.n997 vss 0.150341
R1844 vss.n759 vss.n435 0.14931
R1845 vss.n198 vss.n197 0.145237
R1846 vss.n100 vss.n99 0.145237
R1847 vss.n434 vss.n433 0.145237
R1848 vss.n449 vss.n436 0.139389
R1849 vss.n431 vss.n430 0.133357
R1850 vss.n195 vss.n124 0.133357
R1851 vss.n195 vss.n194 0.133357
R1852 vss.n958 vss.n957 0.133357
R1853 vss.n957 vss.n956 0.133357
R1854 vss.n397 vss.n396 0.133357
R1855 vss.n431 vss.n235 0.133357
R1856 vss.n351 vss 0.126904
R1857 vss vss.n940 0.124938
R1858 vss vss.n199 0.123766
R1859 vss.n757 vss.n435 0.112203
R1860 vss.n1 vss 0.111032
R1861 vss.n759 vss.n758 0.110619
R1862 vss.n687 vss.n686 0.109875
R1863 vss.n689 vss.n688 0.109875
R1864 vss.n746 vss.n644 0.109875
R1865 vss.n737 vss.n736 0.109875
R1866 vss.n572 vss.n571 0.109875
R1867 vss.n597 vss.n596 0.109875
R1868 vss.n500 vss.n499 0.109875
R1869 vss.n787 vss.n786 0.109875
R1870 vss.n752 vss 0.109094
R1871 vss.n349 vss 0.10256
R1872 vss.n510 vss.n451 0.0903438
R1873 vss.n224 vss.n223 0.0860255
R1874 vss.n393 vss.n392 0.0803611
R1875 vss.n750 vss.n749 0.0780862
R1876 vss.n636 vss.n635 0.0780862
R1877 vss.n200 vss 0.0759438
R1878 vss.n450 vss 0.0699444
R1879 vss.n436 vss 0.0699444
R1880 vss.n396 vss.n351 0.0677619
R1881 vss.n994 vss.n993 0.0651358
R1882 vss.n942 vss.n941 0.0651358
R1883 vss.n941 vss 0.0651358
R1884 vss.n421 vss.n420 0.0651358
R1885 vss.n421 vss 0.0651358
R1886 vss.n394 vss.n393 0.0624048
R1887 vss.n3 vss 0.0620278
R1888 vss.n396 vss.n395 0.0576429
R1889 vss.n995 vss 0.0572671
R1890 vss vss.n687 0.0551875
R1891 vss.n688 vss 0.0551875
R1892 vss.n571 vss 0.0551875
R1893 vss vss.n597 0.0551875
R1894 vss vss.n489 0.0551875
R1895 vss.n499 vss 0.0551875
R1896 vss.n223 vss 0.0551875
R1897 vss.n786 vss 0.0551875
R1898 vss vss.n350 0.0524663
R1899 vss.n598 vss 0.0434688
R1900 vss vss.n453 0.0434688
R1901 vss.n350 vss 0.0433241
R1902 vss.n940 vss.n198 0.042429
R1903 vss.n350 vss.n349 0.0417809
R1904 vss.n349 vss.n200 0.0416985
R1905 vss.n747 vss.n642 0.0395625
R1906 vss.n734 vss.n641 0.0354764
R1907 vss.n754 vss.n638 0.034875
R1908 vss vss 0.0346797
R1909 vss.n939 vss.n938 0.0316884
R1910 vss.n736 vss.n735 0.0309688
R1911 vss vss.n724 0.0301875
R1912 vss.n435 vss 0.0297969
R1913 vss.n939 vss.n199 0.0294694
R1914 vss.n758 vss.n450 0.0292698
R1915 vss.n724 vss.n644 0.0255
R1916 vss.n735 vss 0.0247187
R1917 vss.n773 vss.n224 0.0233551
R1918 vss vss.n997 0.0207018
R1919 vss.n489 vss.n451 0.0200312
R1920 vss.n392 vss.n3 0.0188333
R1921 vss.n937 vss.n200 0.0120878
R1922 vss vss.n996 0.00952437
R1923 vss.n995 vss.n994 0.00836871
R1924 vss.n637 vss 0.00513139
R1925 vss.n747 vss 0.00440625
R1926 vss.n635 vss 0.00284375
R1927 vss.n938 vss.n937 0.000993097
R1928 vdd.n600 vdd.n580 5809.41
R1929 vdd.n643 vdd.n600 5809.41
R1930 vdd.n682 vdd.n501 5809.41
R1931 vdd.n501 vdd.n498 5809.41
R1932 vdd.n726 vdd.n691 5809.41
R1933 vdd.n726 vdd.n692 5809.41
R1934 vdd.n729 vdd.n728 5809.41
R1935 vdd.n728 vdd.n483 5809.41
R1936 vdd.n497 vdd.n495 5809.41
R1937 vdd.n684 vdd.n495 5809.41
R1938 vdd.n787 vdd.n39 5809.41
R1939 vdd.n787 vdd.n40 5809.41
R1940 vdd.n815 vdd.n16 5809.41
R1941 vdd.n16 vdd.n13 5809.41
R1942 vdd.n627 vdd.n624 5784.71
R1943 vdd.n628 vdd.n627 5784.71
R1944 vdd.n553 vdd.n487 5784.71
R1945 vdd.n551 vdd.n487 5784.71
R1946 vdd.n713 vdd.n708 5784.71
R1947 vdd.n709 vdd.n708 5784.71
R1948 vdd.n706 vdd.n697 5784.71
R1949 vdd.n706 vdd.n698 5784.71
R1950 vdd.n689 vdd.n489 5784.71
R1951 vdd.n689 vdd.n490 5784.71
R1952 vdd.n70 vdd.n55 5784.71
R1953 vdd.n57 vdd.n55 5784.71
R1954 vdd.n807 vdd.n26 5784.71
R1955 vdd.n809 vdd.n26 5784.71
R1956 vdd.n597 vdd.n585 4912.94
R1957 vdd.n589 vdd.n585 4912.94
R1958 vdd.n597 vdd.n586 4912.94
R1959 vdd.n640 vdd.n603 4912.94
R1960 vdd.n640 vdd.n639 4912.94
R1961 vdd.n639 vdd.n604 4912.94
R1962 vdd.n604 vdd.n603 4912.94
R1963 vdd.n674 vdd.n513 4912.94
R1964 vdd.n674 vdd.n514 4912.94
R1965 vdd.n513 vdd.n509 4912.94
R1966 vdd.n514 vdd.n509 4912.94
R1967 vdd.n506 vdd.n505 4912.94
R1968 vdd.n677 vdd.n505 4912.94
R1969 vdd.n676 vdd.n506 4912.94
R1970 vdd.n677 vdd.n676 4912.94
R1971 vdd.n743 vdd.n469 4912.94
R1972 vdd.n722 vdd.n469 4912.94
R1973 vdd.n743 vdd.n470 4912.94
R1974 vdd.n722 vdd.n470 4912.94
R1975 vdd.n741 vdd.n472 4912.94
R1976 vdd.n720 vdd.n472 4912.94
R1977 vdd.n741 vdd.n473 4912.94
R1978 vdd.n720 vdd.n473 4912.94
R1979 vdd.n796 vdd.n792 4912.94
R1980 vdd.n794 vdd.n792 4912.94
R1981 vdd.n53 vdd.n52 4912.94
R1982 vdd.n76 vdd.n52 4912.94
R1983 vdd.n73 vdd.n53 4912.94
R1984 vdd.n76 vdd.n73 4912.94
R1985 vdd.n794 vdd.n793 4849.41
R1986 vdd.n613 vdd.n612 4207.06
R1987 vdd.n579 vdd.n577 4207.06
R1988 vdd.n646 vdd.n577 4207.06
R1989 vdd.n636 vdd.n613 4207.06
R1990 vdd.n561 vdd.n541 4207.06
R1991 vdd.n541 vdd.n540 4207.06
R1992 vdd.n665 vdd.n536 4207.06
R1993 vdd.n665 vdd.n664 4207.06
R1994 vdd.n747 vdd.n460 4207.06
R1995 vdd.n749 vdd.n460 4207.06
R1996 vdd.n755 vdd.n456 4207.06
R1997 vdd.n456 vdd.n452 4207.06
R1998 vdd.n522 vdd.n519 4207.06
R1999 vdd.n523 vdd.n522 4207.06
R2000 vdd.n667 vdd.n524 4207.06
R2001 vdd.n668 vdd.n667 4207.06
R2002 vdd.n475 vdd.n465 4207.06
R2003 vdd.n475 vdd.n463 4207.06
R2004 vdd.n757 vdd.n450 4207.06
R2005 vdd.n453 vdd.n450 4207.06
R2006 vdd.n791 vdd.n33 4207.06
R2007 vdd.n803 vdd.n791 4207.06
R2008 vdd.n67 vdd.n61 4207.06
R2009 vdd.n61 vdd.n59 4207.06
R2010 vdd.n775 vdd.n80 4207.06
R2011 vdd.n776 vdd.n775 4207.06
R2012 vdd.n624 vdd.n616 4020
R2013 vdd.n628 vdd.n582 4020
R2014 vdd.n553 vdd.n500 4020
R2015 vdd.n551 vdd.n550 4020
R2016 vdd.n713 vdd.n712 4020
R2017 vdd.n710 vdd.n709 4020
R2018 vdd.n697 vdd.n482 4020
R2019 vdd.n700 vdd.n698 4020
R2020 vdd.n510 vdd.n489 4020
R2021 vdd.n494 vdd.n490 4020
R2022 vdd.n70 vdd.n44 4020
R2023 vdd.n57 vdd.n45 4020
R2024 vdd.n807 vdd.n15 4020
R2025 vdd.n810 vdd.n809 4020
R2026 vdd.n616 vdd.n580 3998.82
R2027 vdd.n643 vdd.n582 3998.82
R2028 vdd.n682 vdd.n500 3998.82
R2029 vdd.n550 vdd.n498 3998.82
R2030 vdd.n712 vdd.n691 3998.82
R2031 vdd.n710 vdd.n692 3998.82
R2032 vdd.n729 vdd.n482 3998.82
R2033 vdd.n700 vdd.n483 3998.82
R2034 vdd.n510 vdd.n497 3998.82
R2035 vdd.n684 vdd.n494 3998.82
R2036 vdd.n44 vdd.n39 3998.82
R2037 vdd.n45 vdd.n40 3998.82
R2038 vdd.n815 vdd.n15 3998.82
R2039 vdd.n810 vdd.n13 3998.82
R2040 vdd.n818 vdd.n10 3734.12
R2041 vdd.n612 vdd.n611 3409.41
R2042 vdd.n611 vdd.n579 3409.41
R2043 vdd.n636 vdd.n576 3409.41
R2044 vdd.n646 vdd.n576 3409.41
R2045 vdd.n562 vdd.n561 3409.41
R2046 vdd.n562 vdd.n536 3409.41
R2047 vdd.n540 vdd.n537 3409.41
R2048 vdd.n664 vdd.n537 3409.41
R2049 vdd.n747 vdd.n455 3409.41
R2050 vdd.n755 vdd.n455 3409.41
R2051 vdd.n750 vdd.n749 3409.41
R2052 vdd.n750 vdd.n452 3409.41
R2053 vdd.n519 vdd.n518 3409.41
R2054 vdd.n524 vdd.n518 3409.41
R2055 vdd.n669 vdd.n523 3409.41
R2056 vdd.n669 vdd.n668 3409.41
R2057 vdd.n465 vdd.n449 3409.41
R2058 vdd.n757 vdd.n449 3409.41
R2059 vdd.n733 vdd.n463 3409.41
R2060 vdd.n733 vdd.n453 3409.41
R2061 vdd.n33 vdd.n9 3409.41
R2062 vdd.n818 vdd.n9 3409.41
R2063 vdd.n803 vdd.n802 3409.41
R2064 vdd.n802 vdd.n12 3409.41
R2065 vdd.n67 vdd.n48 3409.41
R2066 vdd.n80 vdd.n48 3409.41
R2067 vdd.n59 vdd.n49 3409.41
R2068 vdd.n776 vdd.n49 3409.41
R2069 vdd.n618 vdd.n616 1789.41
R2070 vdd.n618 vdd.n582 1789.41
R2071 vdd.n433 vdd.n407 1789.41
R2072 vdd.n407 vdd.n403 1789.41
R2073 vdd.n433 vdd.n408 1789.41
R2074 vdd.n408 vdd.n403 1789.41
R2075 vdd.n406 vdd.n400 1789.41
R2076 vdd.n435 vdd.n400 1789.41
R2077 vdd.n406 vdd.n401 1789.41
R2078 vdd.n435 vdd.n401 1789.41
R2079 vdd.n416 vdd.n411 1789.41
R2080 vdd.n425 vdd.n411 1789.41
R2081 vdd.n416 vdd.n412 1789.41
R2082 vdd.n425 vdd.n412 1789.41
R2083 vdd.n418 vdd.n414 1789.41
R2084 vdd.n423 vdd.n418 1789.41
R2085 vdd.n419 vdd.n414 1789.41
R2086 vdd.n423 vdd.n419 1789.41
R2087 vdd.n153 vdd.n141 1789.41
R2088 vdd.n150 vdd.n141 1789.41
R2089 vdd.n153 vdd.n142 1789.41
R2090 vdd.n159 vdd.n136 1789.41
R2091 vdd.n156 vdd.n136 1789.41
R2092 vdd.n159 vdd.n137 1789.41
R2093 vdd.n156 vdd.n137 1789.41
R2094 vdd.n123 vdd.n94 1789.41
R2095 vdd.n123 vdd.n95 1789.41
R2096 vdd.n163 vdd.n87 1789.41
R2097 vdd.n134 vdd.n87 1789.41
R2098 vdd.n116 vdd.n97 1789.41
R2099 vdd.n119 vdd.n97 1789.41
R2100 vdd.n116 vdd.n98 1789.41
R2101 vdd.n119 vdd.n98 1789.41
R2102 vdd.n113 vdd.n102 1789.41
R2103 vdd.n110 vdd.n103 1789.41
R2104 vdd.n113 vdd.n103 1789.41
R2105 vdd.n549 vdd.n500 1789.41
R2106 vdd.n550 vdd.n549 1789.41
R2107 vdd.n712 vdd.n711 1789.41
R2108 vdd.n711 vdd.n710 1789.41
R2109 vdd.n701 vdd.n482 1789.41
R2110 vdd.n701 vdd.n700 1789.41
R2111 vdd.n511 vdd.n510 1789.41
R2112 vdd.n511 vdd.n494 1789.41
R2113 vdd.n782 vdd.n44 1789.41
R2114 vdd.n782 vdd.n45 1789.41
R2115 vdd.n811 vdd.n15 1789.41
R2116 vdd.n811 vdd.n810 1789.41
R2117 vdd.n203 vdd.n188 1789.41
R2118 vdd.n210 vdd.n188 1789.41
R2119 vdd.n203 vdd.n189 1789.41
R2120 vdd.n210 vdd.n189 1789.41
R2121 vdd.n219 vdd.n181 1789.41
R2122 vdd.n200 vdd.n181 1789.41
R2123 vdd.n219 vdd.n182 1789.41
R2124 vdd.n200 vdd.n182 1789.41
R2125 vdd.n331 vdd.n324 1789.41
R2126 vdd.n324 vdd.n322 1789.41
R2127 vdd.n343 vdd.n176 1789.41
R2128 vdd.n345 vdd.n176 1789.41
R2129 vdd.n305 vdd.n286 1789.41
R2130 vdd.n305 vdd.n287 1789.41
R2131 vdd.n319 vdd.n245 1789.41
R2132 vdd.n319 vdd.n246 1789.41
R2133 vdd.n279 vdd.n251 1789.41
R2134 vdd.n308 vdd.n251 1789.41
R2135 vdd.n279 vdd.n252 1789.41
R2136 vdd.n308 vdd.n252 1789.41
R2137 vdd.n271 vdd.n263 1789.41
R2138 vdd.n263 vdd.n258 1789.41
R2139 vdd.n271 vdd.n264 1789.41
R2140 vdd.n264 vdd.n258 1789.41
R2141 vdd.n205 vdd.n191 1789.41
R2142 vdd.n208 vdd.n191 1789.41
R2143 vdd.n205 vdd.n192 1789.41
R2144 vdd.n208 vdd.n192 1789.41
R2145 vdd.n194 vdd.n179 1789.41
R2146 vdd.n199 vdd.n194 1789.41
R2147 vdd.n195 vdd.n179 1789.41
R2148 vdd.n199 vdd.n195 1789.41
R2149 vdd.n323 vdd.n242 1789.41
R2150 vdd.n333 vdd.n242 1789.41
R2151 vdd.n238 vdd.n222 1789.41
R2152 vdd.n238 vdd.n178 1789.41
R2153 vdd.n281 vdd.n254 1789.41
R2154 vdd.n284 vdd.n254 1789.41
R2155 vdd.n281 vdd.n255 1789.41
R2156 vdd.n284 vdd.n255 1789.41
R2157 vdd.n273 vdd.n259 1789.41
R2158 vdd.n276 vdd.n259 1789.41
R2159 vdd.n273 vdd.n260 1789.41
R2160 vdd.n276 vdd.n260 1789.41
R2161 vdd.n389 vdd.n363 1789.41
R2162 vdd.n363 vdd.n359 1789.41
R2163 vdd.n389 vdd.n364 1789.41
R2164 vdd.n364 vdd.n359 1789.41
R2165 vdd.n362 vdd.n356 1789.41
R2166 vdd.n391 vdd.n356 1789.41
R2167 vdd.n362 vdd.n357 1789.41
R2168 vdd.n391 vdd.n357 1789.41
R2169 vdd.n372 vdd.n367 1789.41
R2170 vdd.n381 vdd.n367 1789.41
R2171 vdd.n372 vdd.n368 1789.41
R2172 vdd.n381 vdd.n368 1789.41
R2173 vdd.n374 vdd.n370 1789.41
R2174 vdd.n379 vdd.n374 1789.41
R2175 vdd.n375 vdd.n370 1789.41
R2176 vdd.n379 vdd.n375 1789.41
R2177 vdd.n598 vdd.n584 1534.21
R2178 vdd.n122 vdd.n120 1315.04
R2179 vdd.n89 vdd.n86 1231.76
R2180 vdd.n90 vdd.n89 1231.76
R2181 vdd.n129 vdd.n128 1231.76
R2182 vdd.n128 vdd.n92 1231.76
R2183 vdd.n224 vdd.n223 1231.76
R2184 vdd.n223 vdd.n175 1231.76
R2185 vdd.n326 vdd.n226 1231.76
R2186 vdd.n326 vdd.n325 1231.76
R2187 vdd.n295 vdd.n294 1231.76
R2188 vdd.n294 vdd.n293 1231.76
R2189 vdd.n300 vdd.n289 1231.76
R2190 vdd.n300 vdd.n290 1231.76
R2191 vdd.n234 vdd.n231 1231.76
R2192 vdd.n234 vdd.n233 1231.76
R2193 vdd.n335 vdd.n230 1231.76
R2194 vdd.n335 vdd.n334 1231.76
R2195 vdd.n589 vdd.n588 1189.42
R2196 vdd.n611 vdd.n610 797.648
R2197 vdd.n610 vdd.n576 797.648
R2198 vdd.n563 vdd.n562 797.648
R2199 vdd.n563 vdd.n537 797.648
R2200 vdd.n751 vdd.n455 797.648
R2201 vdd.n751 vdd.n750 797.648
R2202 vdd.n670 vdd.n518 797.648
R2203 vdd.n670 vdd.n669 797.648
R2204 vdd.n734 vdd.n449 797.648
R2205 vdd.n734 vdd.n733 797.648
R2206 vdd.n801 vdd.n9 797.648
R2207 vdd.n802 vdd.n801 797.648
R2208 vdd.n780 vdd.n48 797.648
R2209 vdd.n780 vdd.n49 797.648
R2210 vdd.n129 vdd.n94 557.648
R2211 vdd.n130 vdd.n129 557.648
R2212 vdd.n130 vdd.n86 557.648
R2213 vdd.n163 vdd.n86 557.648
R2214 vdd.n95 vdd.n92 557.648
R2215 vdd.n132 vdd.n92 557.648
R2216 vdd.n132 vdd.n90 557.648
R2217 vdd.n134 vdd.n90 557.648
R2218 vdd.n331 vdd.n226 557.648
R2219 vdd.n341 vdd.n226 557.648
R2220 vdd.n341 vdd.n224 557.648
R2221 vdd.n343 vdd.n224 557.648
R2222 vdd.n325 vdd.n322 557.648
R2223 vdd.n325 vdd.n228 557.648
R2224 vdd.n228 vdd.n175 557.648
R2225 vdd.n345 vdd.n175 557.648
R2226 vdd.n289 vdd.n286 557.648
R2227 vdd.n297 vdd.n289 557.648
R2228 vdd.n297 vdd.n295 557.648
R2229 vdd.n295 vdd.n245 557.648
R2230 vdd.n290 vdd.n287 557.648
R2231 vdd.n291 vdd.n290 557.648
R2232 vdd.n293 vdd.n291 557.648
R2233 vdd.n293 vdd.n246 557.648
R2234 vdd.n323 vdd.n230 557.648
R2235 vdd.n339 vdd.n230 557.648
R2236 vdd.n339 vdd.n231 557.648
R2237 vdd.n231 vdd.n222 557.648
R2238 vdd.n334 vdd.n333 557.648
R2239 vdd.n334 vdd.n229 557.648
R2240 vdd.n233 vdd.n229 557.648
R2241 vdd.n233 vdd.n178 557.648
R2242 vdd vdd.n587 524.352
R2243 vdd.n596 vdd.n587 524.068
R2244 vdd.n5 vdd.n4 486.526
R2245 vdd.n590 vdd 478.745
R2246 vdd.n599 vdd.n598 473.772
R2247 vdd.n596 vdd.n595 473.219
R2248 vdd.n621 vdd.n620 447.06
R2249 vdd.n681 vdd.n680 447.06
R2250 vdd.n725 vdd.n716 447.06
R2251 vdd.n699 vdd.n485 447.06
R2252 vdd.n685 vdd.n493 447.06
R2253 vdd.n786 vdd.n785 447.06
R2254 vdd.n24 vdd.n23 447.06
R2255 vdd.n623 vdd.n614 444.515
R2256 vdd.n555 vdd.n554 444.515
R2257 vdd.n714 vdd.n696 444.515
R2258 vdd.n705 vdd.n704 444.515
R2259 vdd.n688 vdd.n687 444.515
R2260 vdd.n62 vdd.n42 444.515
R2261 vdd.n35 vdd.n27 444.515
R2262 vdd.n623 vdd.n622 428.8
R2263 vdd.n554 vdd.n502 428.8
R2264 vdd.n715 vdd.n714 428.8
R2265 vdd.n704 vdd.n703 428.8
R2266 vdd.n687 vdd.n686 428.8
R2267 vdd.n784 vdd.n42 428.8
R2268 vdd.n27 vdd.n25 428.8
R2269 vdd.n622 vdd.n621 426.541
R2270 vdd.n681 vdd.n502 426.541
R2271 vdd.n716 vdd.n715 426.541
R2272 vdd.n703 vdd.n699 426.541
R2273 vdd.n686 vdd.n685 426.541
R2274 vdd.n785 vdd.n784 426.541
R2275 vdd.n25 vdd.n24 426.541
R2276 vdd.n819 vdd.n8 378.38
R2277 vdd.n635 vdd.n574 363.671
R2278 vdd.n565 vdd.n538 363.671
R2279 vdd.n461 vdd.n459 363.671
R2280 vdd.n474 vdd.n447 363.671
R2281 vdd.n520 vdd.n517 363.671
R2282 vdd.n66 vdd.n50 363.671
R2283 vdd.n34 vdd.n7 363.671
R2284 vdd.n648 vdd.n647 363.295
R2285 vdd.n663 vdd.n662 363.295
R2286 vdd.n717 vdd.n444 363.295
R2287 vdd.n759 vdd.n758 363.295
R2288 vdd.n568 vdd.n567 363.295
R2289 vdd.n773 vdd.n772 363.295
R2290 vdd.n820 vdd.n819 363.295
R2291 vdd.n635 vdd.n634 362.37
R2292 vdd.n556 vdd.n538 362.37
R2293 vdd.n521 vdd.n520 362.37
R2294 vdd.n467 vdd.n461 362.37
R2295 vdd.n476 vdd.n474 362.37
R2296 vdd.n37 vdd.n34 362.37
R2297 vdd.n66 vdd.n65 362.37
R2298 vdd.n647 vdd.n575 361.584
R2299 vdd.n663 vdd.n503 361.584
R2300 vdd.n567 vdd.n534 361.584
R2301 vdd.n718 vdd.n717 361.584
R2302 vdd.n758 vdd.n448 361.584
R2303 vdd.n774 vdd.n773 361.584
R2304 vdd.n645 vdd.n578 349.733
R2305 vdd.n781 vdd.n47 349.733
R2306 vdd.n817 vdd.n11 349.733
R2307 vdd.n638 vdd.n637 341.769
R2308 vdd.n68 vdd.n46 341.769
R2309 vdd.n795 vdd.n29 341.769
R2310 vdd.n789 vdd.n788 304.478
R2311 vdd.n32 vdd.n31 294.932
R2312 vdd.n583 vdd.n581 285.291
R2313 vdd.n75 vdd.n38 285.291
R2314 vdd.n626 vdd.n625 269.361
R2315 vdd.n60 vdd.n56 269.361
R2316 vdd.n790 vdd.n28 269.361
R2317 vdd.n19 vdd.n14 245.827
R2318 vdd.n10 vdd.n8 201.326
R2319 vdd.n622 vdd.n619 190.871
R2320 vdd.n619 vdd.n617 190.871
R2321 vdd.n432 vdd 190.871
R2322 vdd.n409 vdd 190.871
R2323 vdd.n432 vdd.n431 190.871
R2324 vdd.n405 vdd 190.871
R2325 vdd.n436 vdd 190.871
R2326 vdd.n405 vdd.n399 190.871
R2327 vdd.n415 vdd.n410 190.871
R2328 vdd.n415 vdd 190.871
R2329 vdd.n426 vdd 190.871
R2330 vdd.n422 vdd 190.871
R2331 vdd vdd.n421 190.871
R2332 vdd.n421 vdd.n420 190.871
R2333 vdd.n152 vdd.n143 190.871
R2334 vdd.n152 vdd 190.871
R2335 vdd vdd.n151 190.871
R2336 vdd.n158 vdd.n138 190.871
R2337 vdd.n158 vdd 190.871
R2338 vdd vdd.n157 190.871
R2339 vdd.n125 vdd.n124 190.871
R2340 vdd.n124 vdd 190.871
R2341 vdd.n164 vdd.n85 190.871
R2342 vdd vdd.n85 190.871
R2343 vdd.n117 vdd.n100 190.871
R2344 vdd vdd.n117 190.871
R2345 vdd.n118 vdd 190.871
R2346 vdd.n112 vdd 190.871
R2347 vdd vdd.n111 190.871
R2348 vdd.n111 vdd.n108 190.871
R2349 vdd.n548 vdd.n502 190.871
R2350 vdd.n548 vdd.n547 190.871
R2351 vdd.n715 vdd.n695 190.871
R2352 vdd.n695 vdd.n694 190.871
R2353 vdd.n702 vdd.n480 190.871
R2354 vdd.n703 vdd.n702 190.871
R2355 vdd.n529 vdd.n492 190.871
R2356 vdd.n686 vdd.n492 190.871
R2357 vdd.n783 vdd.n43 190.871
R2358 vdd.n784 vdd.n783 190.871
R2359 vdd.n813 vdd.n812 190.871
R2360 vdd.n812 vdd.n25 190.871
R2361 vdd.n202 vdd 190.871
R2362 vdd.n211 vdd 190.871
R2363 vdd.n202 vdd.n187 190.871
R2364 vdd.n218 vdd 190.871
R2365 vdd.n183 vdd 190.871
R2366 vdd.n218 vdd.n217 190.871
R2367 vdd vdd.n330 190.871
R2368 vdd.n330 vdd.n329 190.871
R2369 vdd vdd.n174 190.871
R2370 vdd.n346 vdd.n174 190.871
R2371 vdd.n304 vdd 190.871
R2372 vdd.n304 vdd.n303 190.871
R2373 vdd.n318 vdd 190.871
R2374 vdd.n318 vdd.n317 190.871
R2375 vdd.n278 vdd 190.871
R2376 vdd.n309 vdd 190.871
R2377 vdd.n278 vdd.n250 190.871
R2378 vdd.n270 vdd 190.871
R2379 vdd.n265 vdd 190.871
R2380 vdd.n270 vdd.n269 190.871
R2381 vdd.n206 vdd.n193 190.871
R2382 vdd vdd.n206 190.871
R2383 vdd.n207 vdd 190.871
R2384 vdd.n197 vdd.n196 190.871
R2385 vdd vdd.n197 190.871
R2386 vdd.n198 vdd 190.871
R2387 vdd.n243 vdd.n232 190.871
R2388 vdd vdd.n243 190.871
R2389 vdd.n239 vdd.n237 190.871
R2390 vdd vdd.n239 190.871
R2391 vdd.n282 vdd.n256 190.871
R2392 vdd vdd.n282 190.871
R2393 vdd.n283 vdd 190.871
R2394 vdd.n275 vdd 190.871
R2395 vdd vdd.n274 190.871
R2396 vdd.n274 vdd.n262 190.871
R2397 vdd.n388 vdd 190.871
R2398 vdd.n365 vdd 190.871
R2399 vdd.n388 vdd.n387 190.871
R2400 vdd.n361 vdd 190.871
R2401 vdd.n392 vdd 190.871
R2402 vdd.n361 vdd.n355 190.871
R2403 vdd.n371 vdd.n366 190.871
R2404 vdd.n371 vdd 190.871
R2405 vdd.n382 vdd 190.871
R2406 vdd.n378 vdd 190.871
R2407 vdd vdd.n377 190.871
R2408 vdd.n377 vdd.n376 190.871
R2409 vdd.n430 vdd.n409 190.494
R2410 vdd.n437 vdd.n436 190.494
R2411 vdd.n427 vdd.n426 190.494
R2412 vdd.n422 vdd.n397 190.494
R2413 vdd.n151 vdd.n148 190.494
R2414 vdd.n157 vdd.n139 190.494
R2415 vdd.n118 vdd.n99 190.494
R2416 vdd.n112 vdd.n107 190.494
R2417 vdd.n212 vdd.n211 190.494
R2418 vdd.n216 vdd.n183 190.494
R2419 vdd.n310 vdd.n309 190.494
R2420 vdd.n268 vdd.n265 190.494
R2421 vdd.n207 vdd.n185 190.494
R2422 vdd.n198 vdd.n184 190.494
R2423 vdd.n283 vdd.n249 190.494
R2424 vdd.n275 vdd.n261 190.494
R2425 vdd.n386 vdd.n365 190.494
R2426 vdd.n393 vdd.n392 190.494
R2427 vdd.n383 vdd.n382 190.494
R2428 vdd.n378 vdd.n353 190.494
R2429 vdd.n20 vdd.n10 185
R2430 vdd.n114 vdd.n101 179.118
R2431 vdd.n115 vdd.n96 179.118
R2432 vdd.n120 vdd.n96 179.118
R2433 vdd.n122 vdd.n121 179.118
R2434 vdd.n121 vdd.n93 179.118
R2435 vdd.n131 vdd.n93 179.118
R2436 vdd.n131 vdd.n88 179.118
R2437 vdd.n162 vdd.n88 179.118
R2438 vdd.n162 vdd.n161 179.118
R2439 vdd.n160 vdd.n135 179.118
R2440 vdd.n155 vdd.n135 179.118
R2441 vdd.n154 vdd.n140 179.118
R2442 vdd.n756 vdd.n451 174.868
R2443 vdd.n512 vdd.n496 174.868
R2444 vdd.n110 vdd.n109 173.642
R2445 vdd.n150 vdd.n149 173.642
R2446 vdd.n748 vdd.n464 170.885
R2447 vdd.n675 vdd.n508 170.885
R2448 vdd.n727 vdd.n690 152.239
R2449 vdd.n721 vdd.n486 142.645
R2450 vdd.n666 vdd.n499 142.645
R2451 vdd.n20 vdd.n16 137.326
R2452 vdd.n627 vdd.n626 136.964
R2453 vdd.n60 vdd.n55 136.964
R2454 vdd.n742 vdd.n471 134.68
R2455 vdd.n543 vdd.n488 134.68
R2456 vdd.n165 vdd.n84 131.388
R2457 vdd.n133 vdd.n84 131.388
R2458 vdd.n127 vdd.n126 131.388
R2459 vdd.n127 vdd.n91 131.388
R2460 vdd.n342 vdd.n173 131.388
R2461 vdd.n347 vdd.n173 131.388
R2462 vdd.n327 vdd.n225 131.388
R2463 vdd.n328 vdd.n327 131.388
R2464 vdd.n296 vdd.n247 131.388
R2465 vdd.n316 vdd.n247 131.388
R2466 vdd.n301 vdd.n288 131.388
R2467 vdd.n302 vdd.n301 131.388
R2468 vdd.n236 vdd.n235 131.388
R2469 vdd.n240 vdd.n235 131.388
R2470 vdd.n337 vdd.n336 131.388
R2471 vdd.n336 vdd.n241 131.388
R2472 vdd.n21 vdd.n20 123.334
R2473 vdd.n599 vdd.n583 123.096
R2474 vdd.n788 vdd.n38 123.096
R2475 vdd.n790 vdd.n789 122.733
R2476 vdd.n161 vdd.n160 120.168
R2477 vdd.n115 vdd.n114 117.9
R2478 vdd.n155 vdd.n154 117.9
R2479 vdd.n793 vdd.n17 98.5799
R2480 vdd.n412 vdd 92.5005
R2481 vdd.n417 vdd.n412 92.5005
R2482 vdd.n411 vdd.n410 92.5005
R2483 vdd.n413 vdd.n411 92.5005
R2484 vdd.n401 vdd.n399 92.5005
R2485 vdd.n404 vdd.n401 92.5005
R2486 vdd.n400 vdd 92.5005
R2487 vdd.n402 vdd.n400 92.5005
R2488 vdd.n431 vdd.n408 92.5005
R2489 vdd.n408 vdd.n404 92.5005
R2490 vdd vdd.n407 92.5005
R2491 vdd.n407 vdd.n402 92.5005
R2492 vdd vdd.n419 92.5005
R2493 vdd.n419 vdd.n417 92.5005
R2494 vdd.n420 vdd.n418 92.5005
R2495 vdd.n418 vdd.n413 92.5005
R2496 vdd vdd.n98 92.5005
R2497 vdd.n98 vdd.n96 92.5005
R2498 vdd.n100 vdd.n97 92.5005
R2499 vdd.n97 vdd.n96 92.5005
R2500 vdd.n134 vdd 92.5005
R2501 vdd.n162 vdd.n134 92.5005
R2502 vdd vdd.n132 92.5005
R2503 vdd.n132 vdd.n131 92.5005
R2504 vdd.n95 vdd 92.5005
R2505 vdd.n121 vdd.n95 92.5005
R2506 vdd.n125 vdd.n94 92.5005
R2507 vdd.n121 vdd.n94 92.5005
R2508 vdd.n130 vdd.n83 92.5005
R2509 vdd.n131 vdd.n130 92.5005
R2510 vdd.n164 vdd.n163 92.5005
R2511 vdd.n163 vdd.n162 92.5005
R2512 vdd vdd.n137 92.5005
R2513 vdd.n137 vdd.n135 92.5005
R2514 vdd.n138 vdd.n136 92.5005
R2515 vdd.n136 vdd.n135 92.5005
R2516 vdd vdd.n142 92.5005
R2517 vdd.n143 vdd.n141 92.5005
R2518 vdd.n141 vdd.n140 92.5005
R2519 vdd vdd.n103 92.5005
R2520 vdd.n103 vdd.n101 92.5005
R2521 vdd.n108 vdd.n102 92.5005
R2522 vdd vdd.n255 92.5005
R2523 vdd.n255 vdd.n253 92.5005
R2524 vdd.n256 vdd.n254 92.5005
R2525 vdd.n254 vdd.n253 92.5005
R2526 vdd vdd.n178 92.5005
R2527 vdd.n344 vdd.n178 92.5005
R2528 vdd vdd.n229 92.5005
R2529 vdd.n340 vdd.n229 92.5005
R2530 vdd.n333 vdd 92.5005
R2531 vdd.n333 vdd.n332 92.5005
R2532 vdd.n323 vdd.n232 92.5005
R2533 vdd.n332 vdd.n323 92.5005
R2534 vdd.n339 vdd.n338 92.5005
R2535 vdd.n340 vdd.n339 92.5005
R2536 vdd.n237 vdd.n222 92.5005
R2537 vdd.n344 vdd.n222 92.5005
R2538 vdd vdd.n195 92.5005
R2539 vdd.n195 vdd.n180 92.5005
R2540 vdd.n196 vdd.n194 92.5005
R2541 vdd.n194 vdd.n180 92.5005
R2542 vdd vdd.n192 92.5005
R2543 vdd.n192 vdd.n190 92.5005
R2544 vdd.n193 vdd.n191 92.5005
R2545 vdd.n191 vdd.n190 92.5005
R2546 vdd.n269 vdd.n264 92.5005
R2547 vdd.n264 vdd.n257 92.5005
R2548 vdd vdd.n263 92.5005
R2549 vdd.n263 vdd.n257 92.5005
R2550 vdd.n252 vdd.n250 92.5005
R2551 vdd.n253 vdd.n252 92.5005
R2552 vdd.n251 vdd 92.5005
R2553 vdd.n253 vdd.n251 92.5005
R2554 vdd.n317 vdd.n246 92.5005
R2555 vdd.n246 vdd.n244 92.5005
R2556 vdd.n291 vdd.n248 92.5005
R2557 vdd.n298 vdd.n291 92.5005
R2558 vdd.n303 vdd.n287 92.5005
R2559 vdd.n287 vdd.n285 92.5005
R2560 vdd vdd.n286 92.5005
R2561 vdd.n286 vdd.n285 92.5005
R2562 vdd.n297 vdd 92.5005
R2563 vdd.n298 vdd.n297 92.5005
R2564 vdd vdd.n245 92.5005
R2565 vdd.n245 vdd.n244 92.5005
R2566 vdd.n346 vdd.n345 92.5005
R2567 vdd.n345 vdd.n344 92.5005
R2568 vdd.n228 vdd.n172 92.5005
R2569 vdd.n340 vdd.n228 92.5005
R2570 vdd.n329 vdd.n322 92.5005
R2571 vdd.n332 vdd.n322 92.5005
R2572 vdd.n331 vdd 92.5005
R2573 vdd.n332 vdd.n331 92.5005
R2574 vdd vdd.n341 92.5005
R2575 vdd.n341 vdd.n340 92.5005
R2576 vdd.n343 vdd 92.5005
R2577 vdd.n344 vdd.n343 92.5005
R2578 vdd.n217 vdd.n182 92.5005
R2579 vdd.n182 vdd.n180 92.5005
R2580 vdd vdd.n181 92.5005
R2581 vdd.n181 vdd.n180 92.5005
R2582 vdd.n189 vdd.n187 92.5005
R2583 vdd.n190 vdd.n189 92.5005
R2584 vdd.n188 vdd 92.5005
R2585 vdd.n190 vdd.n188 92.5005
R2586 vdd vdd.n260 92.5005
R2587 vdd.n260 vdd.n257 92.5005
R2588 vdd.n262 vdd.n259 92.5005
R2589 vdd.n259 vdd.n257 92.5005
R2590 vdd.n368 vdd 92.5005
R2591 vdd.n373 vdd.n368 92.5005
R2592 vdd.n367 vdd.n366 92.5005
R2593 vdd.n369 vdd.n367 92.5005
R2594 vdd.n357 vdd.n355 92.5005
R2595 vdd.n360 vdd.n357 92.5005
R2596 vdd.n356 vdd 92.5005
R2597 vdd.n358 vdd.n356 92.5005
R2598 vdd.n387 vdd.n364 92.5005
R2599 vdd.n364 vdd.n360 92.5005
R2600 vdd vdd.n363 92.5005
R2601 vdd.n363 vdd.n358 92.5005
R2602 vdd vdd.n375 92.5005
R2603 vdd.n375 vdd.n373 92.5005
R2604 vdd.n376 vdd.n374 92.5005
R2605 vdd.n374 vdd.n369 92.5005
R2606 vdd.n434 vdd.n402 91.6935
R2607 vdd.n434 vdd.n404 91.6935
R2608 vdd.n424 vdd.n413 91.6935
R2609 vdd.n424 vdd.n417 91.6935
R2610 vdd.n390 vdd.n358 91.6935
R2611 vdd.n390 vdd.n360 91.6935
R2612 vdd.n380 vdd.n369 91.6935
R2613 vdd.n380 vdd.n373 91.6935
R2614 vdd.n272 vdd.n257 89.559
R2615 vdd.n277 vdd.n257 89.559
R2616 vdd.n280 vdd.n253 89.559
R2617 vdd.n307 vdd.n253 89.559
R2618 vdd.n306 vdd.n285 89.559
R2619 vdd.n299 vdd.n285 89.559
R2620 vdd.n299 vdd.n298 89.559
R2621 vdd.n298 vdd.n292 89.559
R2622 vdd.n292 vdd.n244 89.559
R2623 vdd.n320 vdd.n244 89.559
R2624 vdd.n332 vdd.n321 89.559
R2625 vdd.n332 vdd.n227 89.559
R2626 vdd.n340 vdd.n227 89.559
R2627 vdd.n340 vdd.n177 89.559
R2628 vdd.n344 vdd.n177 89.559
R2629 vdd.n344 vdd.n221 89.559
R2630 vdd.n220 vdd.n180 89.559
R2631 vdd.n201 vdd.n180 89.559
R2632 vdd.n204 vdd.n190 89.559
R2633 vdd.n209 vdd.n190 89.559
R2634 vdd.n609 vdd.n608 85.0829
R2635 vdd.n609 vdd.n574 85.0829
R2636 vdd.n564 vdd.n539 85.0829
R2637 vdd.n565 vdd.n564 85.0829
R2638 vdd.n753 vdd.n752 85.0829
R2639 vdd.n752 vdd.n459 85.0829
R2640 vdd.n735 vdd.n447 85.0829
R2641 vdd.n736 vdd.n735 85.0829
R2642 vdd.n671 vdd.n517 85.0829
R2643 vdd.n672 vdd.n671 85.0829
R2644 vdd.n779 vdd.n50 85.0829
R2645 vdd.n779 vdd.n778 85.0829
R2646 vdd.n800 vdd.n7 85.0829
R2647 vdd.n800 vdd.n799 85.0829
R2648 vdd.n149 vdd.n142 79.4196
R2649 vdd.n109 vdd.n102 79.4196
R2650 vdd.n617 vdd.n601 66.7857
R2651 vdd.n547 vdd.n546 66.7857
R2652 vdd.n694 vdd.n457 66.7857
R2653 vdd.n731 vdd.n480 66.7857
R2654 vdd.n530 vdd.n529 66.7857
R2655 vdd.n79 vdd.n43 66.7857
R2656 vdd.n814 vdd.n813 66.7857
R2657 vdd.n814 vdd.n17 66.6358
R2658 vdd.n629 vdd.n615 66.1931
R2659 vdd.n544 vdd.n542 66.1931
R2660 vdd.n693 vdd.n466 66.1931
R2661 vdd.n479 vdd.n478 66.1931
R2662 vdd.n528 vdd.n527 66.1931
R2663 vdd.n72 vdd.n71 66.1931
R2664 vdd.n806 vdd.n18 66.1931
R2665 vdd.n637 vdd.n606 62.6339
R2666 vdd.n69 vdd.n68 62.6339
R2667 vdd.n808 vdd.n29 62.6339
R2668 vdd.n727 vdd.n486 61.5478
R2669 vdd.n666 vdd.n535 61.5478
R2670 vdd.n707 vdd.n471 61.3667
R2671 vdd.n690 vdd.n488 61.3667
R2672 vdd.n645 vdd.n644 60.4616
R2673 vdd.n74 vdd.n47 60.4616
R2674 vdd.n817 vdd.n816 60.4616
R2675 vdd.n307 vdd.n306 60.084
R2676 vdd.n321 vdd.n320 60.084
R2677 vdd.n221 vdd.n220 60.084
R2678 vdd.n126 vdd.n125 59.4829
R2679 vdd.n126 vdd.n83 59.4829
R2680 vdd.n165 vdd.n164 59.4829
R2681 vdd vdd.n91 59.4829
R2682 vdd vdd.n91 59.4829
R2683 vdd.n133 vdd 59.4829
R2684 vdd vdd.n133 59.4829
R2685 vdd vdd.n225 59.4829
R2686 vdd vdd.n225 59.4829
R2687 vdd.n342 vdd 59.4829
R2688 vdd vdd.n342 59.4829
R2689 vdd.n329 vdd.n328 59.4829
R2690 vdd.n328 vdd.n172 59.4829
R2691 vdd.n347 vdd.n346 59.4829
R2692 vdd.n288 vdd 59.4829
R2693 vdd vdd.n288 59.4829
R2694 vdd vdd.n296 59.4829
R2695 vdd.n296 vdd 59.4829
R2696 vdd.n303 vdd.n302 59.4829
R2697 vdd.n302 vdd.n248 59.4829
R2698 vdd.n317 vdd.n316 59.4829
R2699 vdd.n337 vdd.n232 59.4829
R2700 vdd.n338 vdd.n337 59.4829
R2701 vdd.n237 vdd.n236 59.4829
R2702 vdd vdd.n241 59.4829
R2703 vdd.n241 vdd 59.4829
R2704 vdd vdd.n240 59.4829
R2705 vdd.n240 vdd 59.4829
R2706 vdd.n166 vdd.n165 59.1064
R2707 vdd.n348 vdd.n347 59.1064
R2708 vdd.n316 vdd.n315 59.1064
R2709 vdd.n236 vdd.n170 59.1064
R2710 vdd.n280 vdd.n277 58.9504
R2711 vdd.n204 vdd.n201 58.9504
R2712 vdd.n799 vdd.n798 53.6992
R2713 vdd.n608 vdd.n607 52.3937
R2714 vdd.n545 vdd.n539 52.3937
R2715 vdd.n754 vdd.n753 52.3937
R2716 vdd.n736 vdd.n732 52.3937
R2717 vdd.n672 vdd.n516 52.3937
R2718 vdd.n778 vdd.n777 52.3937
R2719 vdd.n630 vdd.n605 51.2005
R2720 vdd.n560 vdd.n507 51.2005
R2721 vdd.n746 vdd.n458 51.2005
R2722 vdd.n738 vdd.n737 51.2005
R2723 vdd.n673 vdd.n515 51.2005
R2724 vdd.n58 vdd.n51 51.2005
R2725 vdd.n804 vdd.n32 48.9418
R2726 vdd.n793 vdd.n14 46.2505
R2727 vdd.n815 vdd.n814 40.0406
R2728 vdd.n20 vdd.n19 39.4632
R2729 vdd vdd.n589 37.0005
R2730 vdd.n597 vdd.n596 37.0005
R2731 vdd.n598 vdd.n597 37.0005
R2732 vdd.n641 vdd.n640 37.0005
R2733 vdd.n640 vdd.n581 37.0005
R2734 vdd.n577 vdd.n575 37.0005
R2735 vdd.n583 vdd.n577 37.0005
R2736 vdd.n634 vdd.n613 37.0005
R2737 vdd.n626 vdd.n613 37.0005
R2738 vdd.n632 vdd.n604 37.0005
R2739 vdd.n625 vdd.n604 37.0005
R2740 vdd.n610 vdd.n609 37.0005
R2741 vdd.n610 vdd.n578 37.0005
R2742 vdd.n720 vdd.n481 37.0005
R2743 vdd.n721 vdd.n720 37.0005
R2744 vdd.n741 vdd.n740 37.0005
R2745 vdd.n742 vdd.n741 37.0005
R2746 vdd.n735 vdd.n734 37.0005
R2747 vdd.n734 vdd.n451 37.0005
R2748 vdd.n450 vdd.n448 37.0005
R2749 vdd.n486 vdd.n450 37.0005
R2750 vdd.n476 vdd.n475 37.0005
R2751 vdd.n475 vdd.n471 37.0005
R2752 vdd.n667 vdd.n534 37.0005
R2753 vdd.n667 vdd.n666 37.0005
R2754 vdd.n522 vdd.n521 37.0005
R2755 vdd.n522 vdd.n488 37.0005
R2756 vdd.n752 vdd.n751 37.0005
R2757 vdd.n751 vdd.n451 37.0005
R2758 vdd.n718 vdd.n456 37.0005
R2759 vdd.n486 vdd.n456 37.0005
R2760 vdd.n467 vdd.n460 37.0005
R2761 vdd.n471 vdd.n460 37.0005
R2762 vdd.n564 vdd.n563 37.0005
R2763 vdd.n563 vdd.n512 37.0005
R2764 vdd.n665 vdd.n503 37.0005
R2765 vdd.n666 vdd.n665 37.0005
R2766 vdd.n556 vdd.n541 37.0005
R2767 vdd.n541 vdd.n488 37.0005
R2768 vdd.n723 vdd.n722 37.0005
R2769 vdd.n722 vdd.n721 37.0005
R2770 vdd.n744 vdd.n743 37.0005
R2771 vdd.n743 vdd.n742 37.0005
R2772 vdd.n678 vdd.n677 37.0005
R2773 vdd.n677 vdd.n499 37.0005
R2774 vdd.n558 vdd.n506 37.0005
R2775 vdd.n543 vdd.n506 37.0005
R2776 vdd.n532 vdd.n514 37.0005
R2777 vdd.n514 vdd.n499 37.0005
R2778 vdd.n525 vdd.n513 37.0005
R2779 vdd.n543 vdd.n513 37.0005
R2780 vdd.n671 vdd.n670 37.0005
R2781 vdd.n670 vdd.n512 37.0005
R2782 vdd.n77 vdd.n76 37.0005
R2783 vdd.n76 vdd.n75 37.0005
R2784 vdd.n63 vdd.n53 37.0005
R2785 vdd.n56 vdd.n53 37.0005
R2786 vdd.n780 vdd.n779 37.0005
R2787 vdd.n781 vdd.n780 37.0005
R2788 vdd.n775 vdd.n774 37.0005
R2789 vdd.n775 vdd.n38 37.0005
R2790 vdd.n65 vdd.n61 37.0005
R2791 vdd.n61 vdd.n60 37.0005
R2792 vdd.n791 vdd.n37 37.0005
R2793 vdd.n791 vdd.n790 37.0005
R2794 vdd.n792 vdd.n30 37.0005
R2795 vdd.n792 vdd.n28 37.0005
R2796 vdd.n801 vdd.n800 37.0005
R2797 vdd.n801 vdd.n11 37.0005
R2798 vdd.n23 vdd.n22 32.7398
R2799 vdd.n748 vdd.n462 31.3172
R2800 vdd.n552 vdd.n508 31.3172
R2801 vdd.n756 vdd.n454 30.2311
R2802 vdd.n683 vdd.n496 30.2311
R2803 vdd.n633 vdd.n614 26.6787
R2804 vdd.n557 vdd.n555 26.6787
R2805 vdd.n696 vdd.n468 26.6787
R2806 vdd.n705 vdd.n477 26.6787
R2807 vdd.n688 vdd.n491 26.6787
R2808 vdd.n64 vdd.n62 26.6787
R2809 vdd.n36 vdd.n35 26.6787
R2810 vdd.n620 vdd.n602 26.63
R2811 vdd.n680 vdd.n679 26.63
R2812 vdd.n725 vdd.n724 26.63
R2813 vdd.n485 vdd.n484 26.63
R2814 vdd.n533 vdd.n493 26.63
R2815 vdd.n786 vdd.n41 26.63
R2816 vdd.n413 vdd.n404 26.5564
R2817 vdd.n369 vdd.n360 26.5564
R2818 vdd.n426 vdd.n425 23.1255
R2819 vdd.n425 vdd.n424 23.1255
R2820 vdd.n416 vdd.n415 23.1255
R2821 vdd.n424 vdd.n416 23.1255
R2822 vdd.n436 vdd.n435 23.1255
R2823 vdd.n435 vdd.n434 23.1255
R2824 vdd.n406 vdd.n405 23.1255
R2825 vdd.n434 vdd.n406 23.1255
R2826 vdd.n409 vdd.n403 23.1255
R2827 vdd.n434 vdd.n403 23.1255
R2828 vdd.n433 vdd.n432 23.1255
R2829 vdd.n434 vdd.n433 23.1255
R2830 vdd.n423 vdd.n422 23.1255
R2831 vdd.n424 vdd.n423 23.1255
R2832 vdd.n421 vdd.n414 23.1255
R2833 vdd.n424 vdd.n414 23.1255
R2834 vdd.n119 vdd.n118 23.1255
R2835 vdd.n120 vdd.n119 23.1255
R2836 vdd.n117 vdd.n116 23.1255
R2837 vdd.n116 vdd.n115 23.1255
R2838 vdd.n128 vdd.n127 23.1255
R2839 vdd.n128 vdd.n93 23.1255
R2840 vdd.n89 vdd.n84 23.1255
R2841 vdd.n89 vdd.n88 23.1255
R2842 vdd.n87 vdd.n85 23.1255
R2843 vdd.n161 vdd.n87 23.1255
R2844 vdd.n124 vdd.n123 23.1255
R2845 vdd.n123 vdd.n122 23.1255
R2846 vdd.n157 vdd.n156 23.1255
R2847 vdd.n156 vdd.n155 23.1255
R2848 vdd.n159 vdd.n158 23.1255
R2849 vdd.n160 vdd.n159 23.1255
R2850 vdd.n151 vdd.n150 23.1255
R2851 vdd.n153 vdd.n152 23.1255
R2852 vdd.n154 vdd.n153 23.1255
R2853 vdd.n113 vdd.n112 23.1255
R2854 vdd.n114 vdd.n113 23.1255
R2855 vdd.n111 vdd.n110 23.1255
R2856 vdd.n284 vdd.n283 23.1255
R2857 vdd.n307 vdd.n284 23.1255
R2858 vdd.n282 vdd.n281 23.1255
R2859 vdd.n281 vdd.n280 23.1255
R2860 vdd.n336 vdd.n335 23.1255
R2861 vdd.n335 vdd.n227 23.1255
R2862 vdd.n235 vdd.n234 23.1255
R2863 vdd.n234 vdd.n177 23.1255
R2864 vdd.n239 vdd.n238 23.1255
R2865 vdd.n238 vdd.n221 23.1255
R2866 vdd.n243 vdd.n242 23.1255
R2867 vdd.n321 vdd.n242 23.1255
R2868 vdd.n199 vdd.n198 23.1255
R2869 vdd.n201 vdd.n199 23.1255
R2870 vdd.n197 vdd.n179 23.1255
R2871 vdd.n220 vdd.n179 23.1255
R2872 vdd.n208 vdd.n207 23.1255
R2873 vdd.n209 vdd.n208 23.1255
R2874 vdd.n206 vdd.n205 23.1255
R2875 vdd.n205 vdd.n204 23.1255
R2876 vdd.n265 vdd.n258 23.1255
R2877 vdd.n277 vdd.n258 23.1255
R2878 vdd.n271 vdd.n270 23.1255
R2879 vdd.n272 vdd.n271 23.1255
R2880 vdd.n309 vdd.n308 23.1255
R2881 vdd.n308 vdd.n307 23.1255
R2882 vdd.n279 vdd.n278 23.1255
R2883 vdd.n280 vdd.n279 23.1255
R2884 vdd.n301 vdd.n300 23.1255
R2885 vdd.n300 vdd.n299 23.1255
R2886 vdd.n294 vdd.n247 23.1255
R2887 vdd.n294 vdd.n292 23.1255
R2888 vdd.n319 vdd.n318 23.1255
R2889 vdd.n320 vdd.n319 23.1255
R2890 vdd.n305 vdd.n304 23.1255
R2891 vdd.n306 vdd.n305 23.1255
R2892 vdd.n327 vdd.n326 23.1255
R2893 vdd.n326 vdd.n227 23.1255
R2894 vdd.n223 vdd.n173 23.1255
R2895 vdd.n223 vdd.n177 23.1255
R2896 vdd.n176 vdd.n174 23.1255
R2897 vdd.n221 vdd.n176 23.1255
R2898 vdd.n330 vdd.n324 23.1255
R2899 vdd.n324 vdd.n321 23.1255
R2900 vdd.n200 vdd.n183 23.1255
R2901 vdd.n201 vdd.n200 23.1255
R2902 vdd.n219 vdd.n218 23.1255
R2903 vdd.n220 vdd.n219 23.1255
R2904 vdd.n211 vdd.n210 23.1255
R2905 vdd.n210 vdd.n209 23.1255
R2906 vdd.n203 vdd.n202 23.1255
R2907 vdd.n204 vdd.n203 23.1255
R2908 vdd.n276 vdd.n275 23.1255
R2909 vdd.n277 vdd.n276 23.1255
R2910 vdd.n274 vdd.n273 23.1255
R2911 vdd.n273 vdd.n272 23.1255
R2912 vdd.n382 vdd.n381 23.1255
R2913 vdd.n381 vdd.n380 23.1255
R2914 vdd.n372 vdd.n371 23.1255
R2915 vdd.n380 vdd.n372 23.1255
R2916 vdd.n392 vdd.n391 23.1255
R2917 vdd.n391 vdd.n390 23.1255
R2918 vdd.n362 vdd.n361 23.1255
R2919 vdd.n390 vdd.n362 23.1255
R2920 vdd.n365 vdd.n359 23.1255
R2921 vdd.n390 vdd.n359 23.1255
R2922 vdd.n389 vdd.n388 23.1255
R2923 vdd.n390 vdd.n389 23.1255
R2924 vdd.n379 vdd.n378 23.1255
R2925 vdd.n380 vdd.n379 23.1255
R2926 vdd.n377 vdd.n370 23.1255
R2927 vdd.n380 vdd.n370 23.1255
R2928 vdd.n798 vdd.n17 19.2575
R2929 vdd.n631 vdd.n630 19.0689
R2930 vdd.n560 vdd.n559 19.0689
R2931 vdd.n746 vdd.n745 19.0689
R2932 vdd.n739 vdd.n738 19.0689
R2933 vdd.n526 vdd.n515 19.0689
R2934 vdd.n58 vdd.n54 19.0689
R2935 vdd.n805 vdd.n804 19.0689
R2936 vdd.n625 vdd.n606 17.7406
R2937 vdd.n69 vdd.n56 17.7406
R2938 vdd.n808 vdd.n28 17.7406
R2939 vdd.n641 vdd.n602 17.4344
R2940 vdd.n679 vdd.n678 17.4344
R2941 vdd.n724 vdd.n723 17.4344
R2942 vdd.n484 vdd.n481 17.4344
R2943 vdd.n533 vdd.n532 17.4344
R2944 vdd.n77 vdd.n41 17.4344
R2945 vdd.n607 vdd.n601 16.8923
R2946 vdd.n530 vdd.n516 16.8923
R2947 vdd.n546 vdd.n545 16.8923
R2948 vdd.n754 vdd.n457 16.8923
R2949 vdd.n732 vdd.n731 16.8923
R2950 vdd.n777 vdd.n79 16.8923
R2951 vdd.n633 vdd.n632 16.6793
R2952 vdd.n558 vdd.n557 16.6793
R2953 vdd.n744 vdd.n468 16.6793
R2954 vdd.n740 vdd.n477 16.6793
R2955 vdd.n525 vdd.n491 16.6793
R2956 vdd.n64 vdd.n63 16.6793
R2957 vdd.n36 vdd.n30 16.6793
R2958 vdd.n627 vdd.n614 14.2313
R2959 vdd.n619 vdd.n618 14.2313
R2960 vdd.n618 vdd.n578 14.2313
R2961 vdd.n620 vdd.n600 14.2313
R2962 vdd.n600 vdd.n599 14.2313
R2963 vdd.n702 vdd.n701 14.2313
R2964 vdd.n701 vdd.n451 14.2313
R2965 vdd.n728 vdd.n485 14.2313
R2966 vdd.n728 vdd.n727 14.2313
R2967 vdd.n706 vdd.n705 14.2313
R2968 vdd.n707 vdd.n706 14.2313
R2969 vdd.n711 vdd.n695 14.2313
R2970 vdd.n711 vdd.n451 14.2313
R2971 vdd.n726 vdd.n725 14.2313
R2972 vdd.n727 vdd.n726 14.2313
R2973 vdd.n708 vdd.n696 14.2313
R2974 vdd.n708 vdd.n707 14.2313
R2975 vdd.n549 vdd.n548 14.2313
R2976 vdd.n549 vdd.n512 14.2313
R2977 vdd.n680 vdd.n501 14.2313
R2978 vdd.n535 vdd.n501 14.2313
R2979 vdd.n555 vdd.n487 14.2313
R2980 vdd.n690 vdd.n487 14.2313
R2981 vdd.n495 vdd.n493 14.2313
R2982 vdd.n535 vdd.n495 14.2313
R2983 vdd.n511 vdd.n492 14.2313
R2984 vdd.n512 vdd.n511 14.2313
R2985 vdd.n689 vdd.n688 14.2313
R2986 vdd.n690 vdd.n689 14.2313
R2987 vdd.n783 vdd.n782 14.2313
R2988 vdd.n782 vdd.n781 14.2313
R2989 vdd.n787 vdd.n786 14.2313
R2990 vdd.n788 vdd.n787 14.2313
R2991 vdd.n62 vdd.n55 14.2313
R2992 vdd.n23 vdd.n16 14.2313
R2993 vdd.n812 vdd.n811 14.2313
R2994 vdd.n811 vdd.n11 14.2313
R2995 vdd.n35 vdd.n26 14.2313
R2996 vdd.n789 vdd.n26 14.2313
R2997 vdd.n22 vdd.n17 12.6319
R2998 vdd.n149 vdd.n140 8.97701
R2999 vdd.n109 vdd.n101 8.97701
R3000 vdd.n742 vdd.n462 8.87055
R3001 vdd.n552 vdd.n543 8.87055
R3002 vdd.n22 vdd.n21 8.1562
R3003 vdd.n638 vdd.n578 7.96544
R3004 vdd.n781 vdd.n46 7.96544
R3005 vdd.n795 vdd.n11 7.96544
R3006 vdd.n630 vdd.n612 7.11588
R3007 vdd.n637 vdd.n612 7.11588
R3008 vdd.n607 vdd.n579 7.11588
R3009 vdd.n645 vdd.n579 7.11588
R3010 vdd.n647 vdd.n646 7.11588
R3011 vdd.n646 vdd.n645 7.11588
R3012 vdd.n636 vdd.n635 7.11588
R3013 vdd.n637 vdd.n636 7.11588
R3014 vdd.n732 vdd.n453 7.11588
R3015 vdd.n756 vdd.n453 7.11588
R3016 vdd.n738 vdd.n463 7.11588
R3017 vdd.n748 vdd.n463 7.11588
R3018 vdd.n474 vdd.n465 7.11588
R3019 vdd.n748 vdd.n465 7.11588
R3020 vdd.n758 vdd.n757 7.11588
R3021 vdd.n757 vdd.n756 7.11588
R3022 vdd.n717 vdd.n452 7.11588
R3023 vdd.n756 vdd.n452 7.11588
R3024 vdd.n749 vdd.n461 7.11588
R3025 vdd.n749 vdd.n748 7.11588
R3026 vdd.n747 vdd.n746 7.11588
R3027 vdd.n748 vdd.n747 7.11588
R3028 vdd.n755 vdd.n754 7.11588
R3029 vdd.n756 vdd.n755 7.11588
R3030 vdd.n664 vdd.n663 7.11588
R3031 vdd.n664 vdd.n496 7.11588
R3032 vdd.n540 vdd.n538 7.11588
R3033 vdd.n540 vdd.n508 7.11588
R3034 vdd.n561 vdd.n560 7.11588
R3035 vdd.n561 vdd.n508 7.11588
R3036 vdd.n545 vdd.n536 7.11588
R3037 vdd.n536 vdd.n496 7.11588
R3038 vdd.n668 vdd.n516 7.11588
R3039 vdd.n668 vdd.n496 7.11588
R3040 vdd.n523 vdd.n515 7.11588
R3041 vdd.n523 vdd.n508 7.11588
R3042 vdd.n520 vdd.n519 7.11588
R3043 vdd.n519 vdd.n508 7.11588
R3044 vdd.n567 vdd.n524 7.11588
R3045 vdd.n524 vdd.n496 7.11588
R3046 vdd.n777 vdd.n776 7.11588
R3047 vdd.n776 vdd.n47 7.11588
R3048 vdd.n59 vdd.n58 7.11588
R3049 vdd.n68 vdd.n59 7.11588
R3050 vdd.n67 vdd.n66 7.11588
R3051 vdd.n68 vdd.n67 7.11588
R3052 vdd.n773 vdd.n80 7.11588
R3053 vdd.n80 vdd.n47 7.11588
R3054 vdd.n798 vdd.n12 7.11588
R3055 vdd.n817 vdd.n12 7.11588
R3056 vdd.n804 vdd.n803 7.11588
R3057 vdd.n803 vdd.n29 7.11588
R3058 vdd.n34 vdd.n33 7.11588
R3059 vdd.n33 vdd.n29 7.11588
R3060 vdd.n819 vdd.n818 7.11588
R3061 vdd.n818 vdd.n817 7.11588
R3062 vdd.n657 vdd 6.74008
R3063 vdd.n824 vdd 6.737
R3064 vdd vdd.n657 6.73352
R3065 vdd.n766 vdd.n1 6.63939
R3066 vdd.n652 vdd.n571 6.63939
R3067 vdd.n590 vdd.n586 5.78175
R3068 vdd.n587 vdd.n585 5.78175
R3069 vdd.n585 vdd.n584 5.78175
R3070 vdd.n615 vdd.n603 5.78175
R3071 vdd.n638 vdd.n603 5.78175
R3072 vdd.n629 vdd.n628 5.78175
R3073 vdd.n628 vdd.n606 5.78175
R3074 vdd.n624 vdd.n623 5.78175
R3075 vdd.n624 vdd.n606 5.78175
R3076 vdd.n621 vdd.n580 5.78175
R3077 vdd.n644 vdd.n580 5.78175
R3078 vdd.n643 vdd.n642 5.78175
R3079 vdd.n644 vdd.n643 5.78175
R3080 vdd.n639 vdd.n605 5.78175
R3081 vdd.n639 vdd.n638 5.78175
R3082 vdd.n699 vdd.n483 5.78175
R3083 vdd.n483 vdd.n454 5.78175
R3084 vdd.n704 vdd.n698 5.78175
R3085 vdd.n698 vdd.n462 5.78175
R3086 vdd.n697 vdd.n478 5.78175
R3087 vdd.n697 vdd.n462 5.78175
R3088 vdd.n730 vdd.n729 5.78175
R3089 vdd.n729 vdd.n454 5.78175
R3090 vdd.n479 vdd.n473 5.78175
R3091 vdd.n473 vdd.n464 5.78175
R3092 vdd.n737 vdd.n472 5.78175
R3093 vdd.n472 vdd.n464 5.78175
R3094 vdd.n470 vdd.n458 5.78175
R3095 vdd.n470 vdd.n464 5.78175
R3096 vdd.n693 vdd.n469 5.78175
R3097 vdd.n469 vdd.n464 5.78175
R3098 vdd.n676 vdd.n507 5.78175
R3099 vdd.n676 vdd.n675 5.78175
R3100 vdd.n544 vdd.n505 5.78175
R3101 vdd.n675 vdd.n505 5.78175
R3102 vdd.n719 vdd.n692 5.78175
R3103 vdd.n692 vdd.n454 5.78175
R3104 vdd.n709 vdd.n466 5.78175
R3105 vdd.n709 vdd.n462 5.78175
R3106 vdd.n714 vdd.n713 5.78175
R3107 vdd.n713 vdd.n462 5.78175
R3108 vdd.n716 vdd.n691 5.78175
R3109 vdd.n691 vdd.n454 5.78175
R3110 vdd.n504 vdd.n498 5.78175
R3111 vdd.n683 vdd.n498 5.78175
R3112 vdd.n551 vdd.n542 5.78175
R3113 vdd.n552 vdd.n551 5.78175
R3114 vdd.n554 vdd.n553 5.78175
R3115 vdd.n553 vdd.n552 5.78175
R3116 vdd.n682 vdd.n681 5.78175
R3117 vdd.n683 vdd.n682 5.78175
R3118 vdd.n531 vdd.n497 5.78175
R3119 vdd.n683 vdd.n497 5.78175
R3120 vdd.n527 vdd.n489 5.78175
R3121 vdd.n552 vdd.n489 5.78175
R3122 vdd.n528 vdd.n509 5.78175
R3123 vdd.n675 vdd.n509 5.78175
R3124 vdd.n685 vdd.n684 5.78175
R3125 vdd.n684 vdd.n683 5.78175
R3126 vdd.n687 vdd.n490 5.78175
R3127 vdd.n552 vdd.n490 5.78175
R3128 vdd.n674 vdd.n673 5.78175
R3129 vdd.n675 vdd.n674 5.78175
R3130 vdd.n785 vdd.n40 5.78175
R3131 vdd.n74 vdd.n40 5.78175
R3132 vdd.n57 vdd.n42 5.78175
R3133 vdd.n69 vdd.n57 5.78175
R3134 vdd.n71 vdd.n70 5.78175
R3135 vdd.n70 vdd.n69 5.78175
R3136 vdd.n78 vdd.n39 5.78175
R3137 vdd.n74 vdd.n39 5.78175
R3138 vdd.n73 vdd.n72 5.78175
R3139 vdd.n73 vdd.n46 5.78175
R3140 vdd.n52 vdd.n51 5.78175
R3141 vdd.n52 vdd.n46 5.78175
R3142 vdd.n816 vdd.n815 5.78175
R3143 vdd.n807 vdd.n806 5.78175
R3144 vdd.n808 vdd.n807 5.78175
R3145 vdd.n794 vdd.n18 5.78175
R3146 vdd.n795 vdd.n794 5.78175
R3147 vdd.n24 vdd.n13 5.78175
R3148 vdd.n816 vdd.n13 5.78175
R3149 vdd.n809 vdd.n27 5.78175
R3150 vdd.n809 vdd.n808 5.78175
R3151 vdd.n797 vdd.n796 5.78175
R3152 vdd.n796 vdd.n795 5.78175
R3153 vdd.n21 vdd.n8 4.93648
R3154 vdd.n595 vdd.n590 4.71629
R3155 vdd.n602 vdd.n575 4.7119
R3156 vdd.n679 vdd.n503 4.7119
R3157 vdd.n534 vdd.n533 4.7119
R3158 vdd.n724 vdd.n718 4.7119
R3159 vdd.n484 vdd.n448 4.7119
R3160 vdd.n774 vdd.n41 4.7119
R3161 vdd.n634 vdd.n633 4.70083
R3162 vdd.n557 vdd.n556 4.70083
R3163 vdd.n521 vdd.n491 4.70083
R3164 vdd.n468 vdd.n467 4.70083
R3165 vdd.n477 vdd.n476 4.70083
R3166 vdd.n37 vdd.n36 4.70083
R3167 vdd.n65 vdd.n64 4.70083
R3168 vdd.n588 vdd.n586 4.37746
R3169 vdd.n644 vdd.n581 3.98297
R3170 vdd.n464 vdd.n451 3.98297
R3171 vdd.n675 vdd.n512 3.98297
R3172 vdd.n75 vdd.n74 3.98297
R3173 vdd.n816 vdd.n14 3.98297
R3174 vdd.n569 vdd 3.52106
R3175 vdd.n762 vdd 3.52106
R3176 vdd.n763 vdd.n443 3.32168
R3177 vdd vdd.n168 3.05185
R3178 vdd.n572 vdd 2.62366
R3179 vdd.n398 vdd 2.3405
R3180 vdd.n398 vdd 2.3405
R3181 vdd.n428 vdd 2.3405
R3182 vdd.n428 vdd 2.3405
R3183 vdd.n146 vdd 2.3405
R3184 vdd.n145 vdd 2.3405
R3185 vdd.n104 vdd 2.3405
R3186 vdd.n106 vdd 2.3405
R3187 vdd.n266 vdd 2.3405
R3188 vdd.n266 vdd 2.3405
R3189 vdd.n312 vdd 2.3405
R3190 vdd.n312 vdd 2.3405
R3191 vdd.n214 vdd 2.3405
R3192 vdd.n214 vdd 2.3405
R3193 vdd.n186 vdd 2.3405
R3194 vdd.n186 vdd 2.3405
R3195 vdd.n354 vdd 2.3405
R3196 vdd.n354 vdd 2.3405
R3197 vdd.n384 vdd 2.3405
R3198 vdd.n384 vdd 2.3405
R3199 vdd.n82 vdd 2.29412
R3200 vdd.n313 vdd 2.29412
R3201 vdd.n171 vdd 2.29412
R3202 vdd.n171 vdd 2.29412
R3203 vdd.n721 vdd.n454 1.99173
R3204 vdd.n683 vdd.n499 1.99173
R3205 vdd.n446 vdd 1.93224
R3206 vdd.n660 vdd 1.93224
R3207 vdd.n107 vdd.n106 1.92169
R3208 vdd.n823 vdd 1.89811
R3209 vdd.n767 vdd 1.89811
R3210 vdd.n438 vdd.n397 1.8605
R3211 vdd.n429 vdd.n427 1.8605
R3212 vdd.n438 vdd.n437 1.8605
R3213 vdd.n430 vdd.n429 1.8605
R3214 vdd.n105 vdd.n99 1.8605
R3215 vdd.n144 vdd.n139 1.8605
R3216 vdd.n148 vdd.n147 1.8605
R3217 vdd.n267 vdd.n261 1.8605
R3218 vdd.n311 vdd.n249 1.8605
R3219 vdd.n215 vdd.n184 1.8605
R3220 vdd.n213 vdd.n185 1.8605
R3221 vdd.n268 vdd.n267 1.8605
R3222 vdd.n311 vdd.n310 1.8605
R3223 vdd.n216 vdd.n215 1.8605
R3224 vdd.n213 vdd.n212 1.8605
R3225 vdd.n394 vdd.n353 1.8605
R3226 vdd.n385 vdd.n383 1.8605
R3227 vdd.n394 vdd.n393 1.8605
R3228 vdd.n386 vdd.n385 1.8605
R3229 vdd.n631 vdd.n629 1.77828
R3230 vdd.n559 vdd.n542 1.77828
R3231 vdd.n745 vdd.n466 1.77828
R3232 vdd.n739 vdd.n478 1.77828
R3233 vdd.n527 vdd.n526 1.77828
R3234 vdd.n71 vdd.n54 1.77828
R3235 vdd.n806 vdd.n805 1.77828
R3236 vdd.n351 vdd.n169 1.76063
R3237 vdd.n440 vdd.n439 1.76063
R3238 vdd.n656 vdd.n655 1.753
R3239 vdd.n654 vdd.n570 1.753
R3240 vdd.n396 vdd.n395 1.75125
R3241 vdd.n827 vdd.n826 1.603
R3242 vdd.n825 vdd.n0 1.603
R3243 vdd.n797 vdd.n32 1.5976
R3244 vdd.n650 vdd 1.43984
R3245 vdd.n588 vdd.n584 1.40064
R3246 vdd.n654 vdd.n653 1.35732
R3247 vdd.n617 vdd.n615 1.3042
R3248 vdd.n547 vdd.n544 1.3042
R3249 vdd.n694 vdd.n693 1.3042
R3250 vdd.n480 vdd.n479 1.3042
R3251 vdd.n529 vdd.n528 1.3042
R3252 vdd.n72 vdd.n43 1.3042
R3253 vdd.n813 vdd.n18 1.3042
R3254 vdd.n352 vdd.n351 1.28995
R3255 vdd.n608 vdd.n605 1.19372
R3256 vdd.n539 vdd.n507 1.19372
R3257 vdd.n753 vdd.n458 1.19372
R3258 vdd.n737 vdd.n736 1.19372
R3259 vdd.n673 vdd.n672 1.19372
R3260 vdd.n778 vdd.n51 1.19372
R3261 vdd.n799 vdd.n797 1.19372
R3262 vdd.n395 vdd.n352 1.06531
R3263 vdd.n573 vdd 1.06379
R3264 vdd.n439 vdd.n438 1.06168
R3265 vdd.n395 vdd.n394 1.06168
R3266 vdd.n439 vdd.n81 1.05594
R3267 vdd.n770 vdd 1.04172
R3268 vdd.n6 vdd 1.04172
R3269 vdd.n441 vdd.n81 0.974078
R3270 vdd.n764 vdd.n442 0.918935
R3271 vdd.n761 vdd 0.890303
R3272 vdd.n566 vdd 0.890303
R3273 vdd.n441 vdd.n440 0.855704
R3274 vdd.n591 vdd 0.85529
R3275 vdd.n768 vdd 0.854351
R3276 vdd.n822 vdd 0.854351
R3277 vdd.n765 vdd.n764 0.781762
R3278 vdd.n571 vdd 0.768852
R3279 vdd.n167 vdd.n166 0.715885
R3280 vdd.n349 vdd.n170 0.715885
R3281 vdd.n315 vdd.n314 0.715885
R3282 vdd.n349 vdd.n348 0.715885
R3283 vdd.n824 vdd 0.69425
R3284 vdd.n766 vdd 0.69425
R3285 vdd.n651 vdd.n650 0.619997
R3286 vdd.n573 vdd.n572 0.619997
R3287 vdd.n765 vdd 0.559955
R3288 vdd.n446 vdd.n445 0.518921
R3289 vdd.n762 vdd.n761 0.518921
R3290 vdd.n569 vdd.n566 0.518921
R3291 vdd.n660 vdd.n659 0.518921
R3292 vdd.n443 vdd 0.505434
R3293 vdd.n658 vdd 0.505434
R3294 vdd.n770 vdd.n769 0.497975
R3295 vdd.n768 vdd.n767 0.497975
R3296 vdd.n823 vdd.n822 0.497975
R3297 vdd.n655 vdd.n0 0.479286
R3298 vdd.n763 vdd 0.467672
R3299 vdd.n657 vdd 0.467461
R3300 vdd.n168 vdd 0.464224
R3301 vdd.n764 vdd.n763 0.426664
R3302 vdd.n314 vdd 0.413
R3303 vdd.n350 vdd.n349 0.410656
R3304 vdd.n648 vdd.n574 0.376971
R3305 vdd.n431 vdd.n430 0.376971
R3306 vdd.n437 vdd.n399 0.376971
R3307 vdd.n427 vdd.n410 0.376971
R3308 vdd.n420 vdd.n397 0.376971
R3309 vdd.n148 vdd.n143 0.376971
R3310 vdd.n139 vdd.n138 0.376971
R3311 vdd.n166 vdd.n83 0.376971
R3312 vdd.n100 vdd.n99 0.376971
R3313 vdd.n108 vdd.n107 0.376971
R3314 vdd.n662 vdd.n565 0.376971
R3315 vdd.n459 vdd.n444 0.376971
R3316 vdd.n759 vdd.n447 0.376971
R3317 vdd.n568 vdd.n517 0.376971
R3318 vdd.n772 vdd.n50 0.376971
R3319 vdd.n820 vdd.n7 0.376971
R3320 vdd.n212 vdd.n187 0.376971
R3321 vdd.n217 vdd.n216 0.376971
R3322 vdd.n348 vdd.n172 0.376971
R3323 vdd.n315 vdd.n248 0.376971
R3324 vdd.n310 vdd.n250 0.376971
R3325 vdd.n269 vdd.n268 0.376971
R3326 vdd.n193 vdd.n185 0.376971
R3327 vdd.n196 vdd.n184 0.376971
R3328 vdd.n338 vdd.n170 0.376971
R3329 vdd.n256 vdd.n249 0.376971
R3330 vdd.n262 vdd.n261 0.376971
R3331 vdd.n387 vdd.n386 0.376971
R3332 vdd.n393 vdd.n355 0.376971
R3333 vdd.n383 vdd.n366 0.376971
R3334 vdd.n376 vdd.n353 0.376971
R3335 vdd.n652 vdd 0.376726
R3336 vdd.n314 vdd.n313 0.360656
R3337 vdd.n349 vdd.n171 0.360656
R3338 vdd.n591 vdd 0.349949
R3339 vdd.n593 vdd 0.344944
R3340 vdd.n442 vdd.n441 0.34097
R3341 vdd.n632 vdd.n631 0.307571
R3342 vdd.n559 vdd.n558 0.307571
R3343 vdd.n745 vdd.n744 0.307571
R3344 vdd.n740 vdd.n739 0.307571
R3345 vdd.n526 vdd.n525 0.307571
R3346 vdd.n63 vdd.n54 0.307571
R3347 vdd.n805 vdd.n30 0.307571
R3348 vdd.n651 vdd 0.304352
R3349 vdd.n595 vdd.n594 0.291125
R3350 vdd.n593 vdd.n592 0.277007
R3351 vdd.n1 vdd 0.27355
R3352 vdd.n594 vdd.n591 0.2731
R3353 vdd.n2 vdd 0.272663
R3354 vdd.n440 vdd.n396 0.264604
R3355 vdd.n396 vdd.n169 0.263158
R3356 vdd.n445 vdd 0.254776
R3357 vdd.n659 vdd 0.254776
R3358 vdd.n6 vdd.n5 0.249237
R3359 vdd.n5 vdd.n3 0.249237
R3360 vdd.n769 vdd 0.244503
R3361 vdd.n3 vdd 0.244503
R3362 vdd.n352 vdd.n81 0.233429
R3363 vdd.n168 vdd.n167 0.22821
R3364 vdd.n167 vdd.n82 0.201986
R3365 vdd.n642 vdd.n641 0.178728
R3366 vdd.n678 vdd.n504 0.178728
R3367 vdd.n723 vdd.n719 0.178728
R3368 vdd.n730 vdd.n481 0.178728
R3369 vdd.n532 vdd.n531 0.178728
R3370 vdd.n78 vdd.n77 0.178728
R3371 vdd.n215 vdd 0.166125
R3372 vdd.n429 vdd 0.164562
R3373 vdd.n311 vdd 0.164562
R3374 vdd vdd.n213 0.164562
R3375 vdd.n385 vdd 0.164562
R3376 vdd vdd.n824 0.148
R3377 vdd.n761 vdd.n760 0.147704
R3378 vdd.n661 vdd.n566 0.147704
R3379 vdd.n760 vdd.n446 0.146059
R3380 vdd.n661 vdd.n660 0.146059
R3381 vdd.n649 vdd.n648 0.133357
R3382 vdd.n760 vdd.n444 0.133357
R3383 vdd.n760 vdd.n759 0.133357
R3384 vdd.n661 vdd.n568 0.133357
R3385 vdd.n662 vdd.n661 0.133357
R3386 vdd.n772 vdd.n771 0.133357
R3387 vdd.n821 vdd.n820 0.133357
R3388 vdd.n445 vdd.n443 0.131257
R3389 vdd.n659 vdd.n658 0.131257
R3390 vdd.n763 vdd.n762 0.131257
R3391 vdd.n657 vdd.n569 0.129612
R3392 vdd.n592 vdd 0.113524
R3393 vdd.n649 vdd.n573 0.110181
R3394 vdd.n438 vdd.n398 0.109875
R3395 vdd.n429 vdd.n428 0.109875
R3396 vdd.n267 vdd.n266 0.109875
R3397 vdd.n312 vdd.n311 0.109875
R3398 vdd.n215 vdd.n214 0.109875
R3399 vdd.n213 vdd.n186 0.109875
R3400 vdd.n394 vdd.n354 0.109875
R3401 vdd.n385 vdd.n384 0.109875
R3402 vdd.n650 vdd.n649 0.108956
R3403 vdd.n657 vdd 0.100037
R3404 vdd.n652 vdd.n651 0.0979265
R3405 vdd.n642 vdd.n601 0.0977152
R3406 vdd.n546 vdd.n504 0.0977152
R3407 vdd.n719 vdd.n457 0.0977152
R3408 vdd.n731 vdd.n730 0.0977152
R3409 vdd.n531 vdd.n530 0.0977152
R3410 vdd.n79 vdd.n78 0.0977152
R3411 vdd.n572 vdd.n571 0.096701
R3412 vdd.n144 vdd 0.0931573
R3413 vdd vdd.n105 0.0922832
R3414 vdd.n147 vdd 0.0922832
R3415 vdd.n592 vdd 0.0847634
R3416 vdd.n771 vdd.n768 0.079844
R3417 vdd.n822 vdd.n821 0.079844
R3418 vdd.n771 vdd.n770 0.0789574
R3419 vdd.n821 vdd.n6 0.0789574
R3420 vdd.n351 vdd.n350 0.0780862
R3421 vdd.n3 vdd.n2 0.0709787
R3422 vdd.n824 vdd.n823 0.0709787
R3423 vdd.n767 vdd.n766 0.0709787
R3424 vdd.n769 vdd.n1 0.0700922
R3425 vdd.n653 vdd 0.0630773
R3426 vdd.n105 vdd.n104 0.0616888
R3427 vdd.n145 vdd.n144 0.0616888
R3428 vdd.n147 vdd.n146 0.0616888
R3429 vdd.n571 vdd.n442 0.0572867
R3430 vdd vdd.n398 0.0551875
R3431 vdd.n428 vdd 0.0551875
R3432 vdd.n266 vdd 0.0551875
R3433 vdd vdd.n312 0.0551875
R3434 vdd.n214 vdd 0.0551875
R3435 vdd.n186 vdd 0.0551875
R3436 vdd vdd.n354 0.0551875
R3437 vdd.n384 vdd 0.0551875
R3438 vdd.n825 vdd 0.0545625
R3439 vdd.n313 vdd 0.0512812
R3440 vdd vdd.n171 0.0512812
R3441 vdd.n653 vdd.n652 0.045162
R3442 vdd.n655 vdd.n654 0.0388531
R3443 vdd.n826 vdd.n1 0.0351875
R3444 vdd vdd.n656 0.0334335
R3445 vdd.n570 vdd.n443 0.0315396
R3446 vdd.n106 vdd 0.0310944
R3447 vdd.n104 vdd 0.0310944
R3448 vdd vdd.n145 0.0310944
R3449 vdd.n146 vdd 0.0310944
R3450 vdd.n766 vdd.n765 0.0298951
R3451 vdd vdd.n82 0.0289091
R3452 vdd.n2 vdd 0.0265417
R3453 vdd.n827 vdd.n0 0.0256039
R3454 vdd.n658 vdd 0.0140031
R3455 vdd.n826 vdd.n825 0.008
R3456 vdd.n658 vdd 0.00744444
R3457 vdd.n169 vdd 0.00538077
R3458 vdd.n594 vdd.n593 0.00440625
R3459 vdd vdd.n827 0.00308012
R3460 vdd.n350 vdd 0.00284375
R3461 vdd.n656 vdd.n570 0.00113131
R3462 vref.n0 vref 2.51601
R3463 vref.n0 vref 2.11902
R3464 vref vref.n1 0.552397
R3465 vref.n1 vref 0.334205
R3466 vref.n1 vref 0.311326
R3467 vref vref.n0 0.188289
R3468 vref.n1 vref 0.0931339
R3469 vref.n1 vref 0.00686574
R3470 comp_p_1/latch_left.n0 comp_p_1/latch_left.t3 114.778
R3471 comp_p_1/latch_left.n0 comp_p_1/latch_left.t2 106.572
R3472 comp_p_1/latch_left.n1 comp_p_1/latch_left.t0 95.1712
R3473 comp_p_1/latch_left.n2 comp_p_1/latch_left.t1 22.0141
R3474 comp_p_1/latch_left.n1 comp_p_1/latch_left.n0 1.72733
R3475 comp_p_1/latch_left comp_p_1/latch_left.n2 0.717514
R3476 comp_p_1/latch_left.n2 comp_p_1/latch_left.n1 0.599169
R3477 d0.n0 d0.t1 556.78
R3478 d0.t1 d0 547.24
R3479 d0 d0.t0 372.113
R3480 d0.n0 d0 9.54008
R3481 d0 d0.n2 4.54809
R3482 d0.n2 d0 4.43618
R3483 d0.n3 d0 0.719145
R3484 d0.n1 d0.n0 0.253625
R3485 d0 d0.n3 0.199411
R3486 d0 d0 0.063
R3487 d0.n2 d0 0.0443144
R3488 d0.n3 d0 0.0262742
R3489 d0 d0 0.0262732
R3490 d0.n1 d0 0.013
R3491 d0.n3 d0 0.00763393
R3492 d0 d0.n1 0.00565464
R3493 vin.n20 vin.t26 899.324
R3494 vin.n38 vin.t22 899.324
R3495 vin.n31 vin.t14 899.324
R3496 vin.n25 vin.t2 899.324
R3497 vin.n2 vin.t6 899.324
R3498 vin.n7 vin.t10 899.324
R3499 vin.n13 vin.t18 899.324
R3500 vin.n21 vin.t26 898.659
R3501 vin.n39 vin.t22 898.659
R3502 vin.n32 vin.t14 898.659
R3503 vin.n26 vin.t2 898.659
R3504 vin.n3 vin.t6 898.659
R3505 vin.n8 vin.t10 898.659
R3506 vin.n14 vin.t18 898.659
R3507 vin.t23 vin.n38 898.442
R3508 vin.t3 vin.n25 898.442
R3509 vin.t7 vin.n2 898.442
R3510 vin.t19 vin.n13 898.442
R3511 vin.t27 vin.n20 898.442
R3512 vin.t15 vin.n31 898.442
R3513 vin.t11 vin.n7 898.442
R3514 vin.n21 vin.t27 897.754
R3515 vin.n39 vin.t23 897.754
R3516 vin.n32 vin.t15 897.754
R3517 vin.n26 vin.t3 897.754
R3518 vin.n3 vin.t7 897.754
R3519 vin.n8 vin.t11 897.754
R3520 vin.n14 vin.t19 897.754
R3521 vin.n18 vin.t24 895.625
R3522 vin.n36 vin.t20 895.625
R3523 vin.n29 vin.t12 895.625
R3524 vin.n23 vin.t0 895.625
R3525 vin.n0 vin.t4 895.625
R3526 vin.n5 vin.t8 895.625
R3527 vin.n11 vin.t16 895.625
R3528 vin.n18 vin.t25 894.172
R3529 vin.n36 vin.t21 894.172
R3530 vin.n29 vin.t13 894.172
R3531 vin.n23 vin.t1 894.172
R3532 vin.n0 vin.t5 894.172
R3533 vin.n5 vin.t9 894.172
R3534 vin.n11 vin.t17 894.172
R3535 vin.n19 vin.n18 6.30807
R3536 vin.n37 vin.n36 6.30807
R3537 vin.n30 vin.n29 6.30807
R3538 vin.n24 vin.n23 6.30807
R3539 vin.n1 vin.n0 6.30807
R3540 vin.n6 vin.n5 6.30807
R3541 vin.n12 vin.n11 6.30807
R3542 vin.n20 vin.n19 5.39021
R3543 vin.n38 vin.n37 5.39021
R3544 vin.n31 vin.n30 5.39021
R3545 vin.n25 vin.n24 5.39021
R3546 vin.n2 vin.n1 5.39021
R3547 vin.n7 vin.n6 5.39021
R3548 vin.n13 vin.n12 5.39021
R3549 vin.n22 vin.n21 5.38653
R3550 vin.n40 vin.n39 5.38653
R3551 vin.n33 vin.n32 5.38653
R3552 vin.n27 vin.n26 5.38653
R3553 vin.n4 vin.n3 5.38653
R3554 vin.n9 vin.n8 5.38653
R3555 vin.n15 vin.n14 5.38653
R3556 vin.n44 vin.n43 5.20469
R3557 vin.n22 vin.n19 5.11108
R3558 vin.n40 vin.n37 5.11108
R3559 vin.n33 vin.n30 5.11108
R3560 vin.n27 vin.n24 5.11108
R3561 vin.n4 vin.n1 5.11108
R3562 vin.n9 vin.n6 5.11108
R3563 vin.n15 vin.n12 5.11108
R3564 vin.n35 vin.n28 4.57467
R3565 vin.n10 vin 4.13219
R3566 vin.n35 vin.n34 3.68222
R3567 vin.n42 vin.n41 3.10272
R3568 vin.n16 vin 2.68025
R3569 vin.n10 vin 2.66582
R3570 vin.n43 vin.n42 2.43775
R3571 vin.n43 vin 1.54614
R3572 vin vin.n16 1.12357
R3573 vin vin.n22 0.870692
R3574 vin vin.n4 0.870692
R3575 vin vin.n9 0.870692
R3576 vin vin.n15 0.870692
R3577 vin.n34 vin.n33 0.837038
R3578 vin.n41 vin.n40 0.726462
R3579 vin.n16 vin.n10 0.70492
R3580 vin.n28 vin.n27 0.668769
R3581 vin.n42 vin.n35 0.533734
R3582 vin.n17 vin 0.468179
R3583 vin vin.n45 0.371278
R3584 vin.n45 vin 0.332981
R3585 vin.n17 vin 0.23608
R3586 vin.n45 vin 0.20608
R3587 vin.n17 vin 0.146164
R3588 vin.n41 vin 0.0482941
R3589 vin.n44 vin.n17 0.0422977
R3590 vin.n45 vin.n44 0.0422977
R3591 vin.n28 vin 0.0391905
R3592 vin.n34 vin 0.0341538
R3593 comp_p_0/out_left.n1 comp_p_0/out_left.t2 145.612
R3594 comp_p_0/out_left.n2 comp_p_0/out_left.t0 143.417
R3595 comp_p_0/out_left.n0 comp_p_0/out_left.t1 29.4286
R3596 comp_p_0/out_left comp_p_0/out_left.n3 11.6041
R3597 comp_p_0/out_left.n3 comp_p_0/out_left.n2 4.33076
R3598 comp_p_0/out_left.n1 comp_p_0/out_left.n0 2.12634
R3599 comp_p_0/out_left.n2 comp_p_0/out_left.n1 2.04428
R3600 comp_p_0/out_left.n3 comp_p_0/out_left.n0 0.00290385
R3601 d1.n0 d1.t1 556.78
R3602 d1.t1 d1 547.24
R3603 d1 d1.t0 372.113
R3604 d1.n1 d1 20.4931
R3605 d1.n0 d1 9.54008
R3606 d1 d1.n1 3.45602
R3607 d1.n2 d1 1.7016
R3608 d1.n1 d1 1.38807
R3609 d1 d1.n2 0.538602
R3610 d1 d1.n0 0.266125
R3611 d1 d1 0.063
R3612 d1.n2 d1 0.0217258
R3613 d1.n2 d1 0.00721429
R3614 comp_p_2/latch_left.n0 comp_p_2/latch_left.t3 114.778
R3615 comp_p_2/latch_left.n0 comp_p_2/latch_left.t2 106.572
R3616 comp_p_2/latch_left.n1 comp_p_2/latch_left.t0 95.1712
R3617 comp_p_2/latch_left.n2 comp_p_2/latch_left.t1 22.0141
R3618 comp_p_2/latch_left.n1 comp_p_2/latch_left.n0 1.72733
R3619 comp_p_2/latch_left comp_p_2/latch_left.n2 0.717514
R3620 comp_p_2/latch_left.n2 comp_p_2/latch_left.n1 0.599169
R3621 d2.n0 d2.t1 556.78
R3622 d2.t1 d2 547.24
R3623 d2 d2.t0 372.113
R3624 d2.n2 d2 18.5756
R3625 d2.n0 d2 9.54008
R3626 d2.n4 d2 2.94937
R3627 d2.n2 d2 1.06075
R3628 d2.n3 d2.n2 0.853
R3629 d2 d2.n4 0.464536
R3630 d2.n1 d2.n0 0.25675
R3631 d2.n4 d2 0.0929839
R3632 d2 d2 0.063
R3633 d2 d2 0.0329675
R3634 d2.n1 d2 0.009875
R3635 d2.n4 d2.n3 0.00777665
R3636 d2.n3 d2 0.00777665
R3637 d2 d2.n1 0.00537013
R3638 comp_p_3/latch_left.n0 comp_p_3/latch_left.t3 114.778
R3639 comp_p_3/latch_left.n0 comp_p_3/latch_left.t2 106.572
R3640 comp_p_3/latch_left.n1 comp_p_3/latch_left.t0 95.1712
R3641 comp_p_3/latch_left.n2 comp_p_3/latch_left.t1 22.0141
R3642 comp_p_3/latch_left.n1 comp_p_3/latch_left.n0 1.72733
R3643 comp_p_3/latch_left comp_p_3/latch_left.n2 0.717514
R3644 comp_p_3/latch_left.n2 comp_p_3/latch_left.n1 0.599169
R3645 comp_p_3/latch_right.n1 comp_p_3/latch_right.t3 114.778
R3646 comp_p_3/latch_right.n1 comp_p_3/latch_right.t2 106.572
R3647 comp_p_3/latch_right.n2 comp_p_3/latch_right.t0 94.6192
R3648 comp_p_3/latch_right.n0 comp_p_3/latch_right.t1 22.0141
R3649 comp_p_3/latch_right.n2 comp_p_3/latch_right.n0 2.37533
R3650 comp_p_3/latch_right.n3 comp_p_3/latch_right.n1 1.43373
R3651 comp_p_3/latch_right.n4 comp_p_3/latch_right.n3 1.11841
R3652 comp_p_3/latch_right.n3 comp_p_3/latch_right.n2 1.06963
R3653 comp_p_3/latch_right comp_p_3/latch_right.n4 0.608139
R3654 comp_p_3/latch_right.n4 comp_p_3/latch_right.n0 0.00530769
R3655 comp_p_3/out_left.n1 comp_p_3/out_left.t2 145.612
R3656 comp_p_3/out_left.n2 comp_p_3/out_left.t0 143.417
R3657 comp_p_3/out_left.n0 comp_p_3/out_left.t1 29.4286
R3658 comp_p_3/out_left comp_p_3/out_left.n3 11.6041
R3659 comp_p_3/out_left.n3 comp_p_3/out_left.n2 4.33076
R3660 comp_p_3/out_left.n1 comp_p_3/out_left.n0 2.12634
R3661 comp_p_3/out_left.n2 comp_p_3/out_left.n1 2.04428
R3662 comp_p_3/out_left.n3 comp_p_3/out_left.n0 0.00290385
R3663 d3.n0 d3.t1 556.78
R3664 d3.t1 d3 547.24
R3665 d3 d3.t0 372.113
R3666 d3.n1 d3 10.0074
R3667 d3.n0 d3 9.54008
R3668 d3.n3 d3 3.8636
R3669 d3.n2 d3.n1 1.978
R3670 d3 d3.n3 1.07938
R3671 d3.n1 d3 0.589103
R3672 d3 d3.n0 0.266125
R3673 d3.n3 d3 0.0975323
R3674 d3 d3 0.063
R3675 d3.n3 d3.n2 0.0223063
R3676 d3.n2 d3 0.00579279
R3677 comp_p_4/latch_left.n0 comp_p_4/latch_left.t3 114.778
R3678 comp_p_4/latch_left.n0 comp_p_4/latch_left.t2 106.572
R3679 comp_p_4/latch_left.n1 comp_p_4/latch_left.t0 95.1712
R3680 comp_p_4/latch_left.n2 comp_p_4/latch_left.t1 22.0141
R3681 comp_p_4/latch_left.n1 comp_p_4/latch_left.n0 1.72733
R3682 comp_p_4/latch_left comp_p_4/latch_left.n2 0.717514
R3683 comp_p_4/latch_left.n2 comp_p_4/latch_left.n1 0.599169
R3684 comp_p_4/out_left.n1 comp_p_4/out_left.t2 145.612
R3685 comp_p_4/out_left.n2 comp_p_4/out_left.t0 143.417
R3686 comp_p_4/out_left.n0 comp_p_4/out_left.t1 29.4286
R3687 comp_p_4/out_left comp_p_4/out_left.n3 11.6041
R3688 comp_p_4/out_left.n3 comp_p_4/out_left.n2 4.33076
R3689 comp_p_4/out_left.n1 comp_p_4/out_left.n0 2.12634
R3690 comp_p_4/out_left.n2 comp_p_4/out_left.n1 2.04428
R3691 comp_p_4/out_left.n3 comp_p_4/out_left.n0 0.00290385
R3692 d4.n0 d4.t1 556.78
R3693 d4.t1 d4 547.24
R3694 d4 d4.t0 372.113
R3695 d4.n1 d4 24.2927
R3696 d4.n0 d4 9.54008
R3697 d4.n2 d4 5.15685
R3698 d4.n1 d4 1.81119
R3699 d4 d4.n2 1.15048
R3700 d4 d4.n1 1.14663
R3701 d4 d4.n0 0.266125
R3702 d4 d4 0.063
R3703 d4.n2 d4 0.00656452
R3704 d4.n2 d4 0.00185252
R3705 comp_p_5/latch_left.n0 comp_p_5/latch_left.t3 114.778
R3706 comp_p_5/latch_left.n0 comp_p_5/latch_left.t2 106.572
R3707 comp_p_5/latch_left.n1 comp_p_5/latch_left.t0 95.1712
R3708 comp_p_5/latch_left.n2 comp_p_5/latch_left.t1 22.0141
R3709 comp_p_5/latch_left.n1 comp_p_5/latch_left.n0 1.72733
R3710 comp_p_5/latch_left comp_p_5/latch_left.n2 0.717514
R3711 comp_p_5/latch_left.n2 comp_p_5/latch_left.n1 0.599169
R3712 d5.n0 d5.t1 556.78
R3713 d5.t1 d5 547.24
R3714 d5 d5.t0 372.113
R3715 d5.n0 d5 9.54008
R3716 d5 d5.n1 3.01518
R3717 d5.n1 d5 2.80934
R3718 d5.n1 d5 0.322375
R3719 d5 d5.n0 0.266125
R3720 d5 d5 0.063
R3721 comp_p_6/latch_left.n0 comp_p_6/latch_left.t3 114.778
R3722 comp_p_6/latch_left.n0 comp_p_6/latch_left.t2 106.572
R3723 comp_p_6/latch_left.n1 comp_p_6/latch_left.t0 95.1712
R3724 comp_p_6/latch_left.n2 comp_p_6/latch_left.t1 22.0141
R3725 comp_p_6/latch_left.n1 comp_p_6/latch_left.n0 1.72733
R3726 comp_p_6/latch_left comp_p_6/latch_left.n2 0.717514
R3727 comp_p_6/latch_left.n2 comp_p_6/latch_left.n1 0.599169
R3728 comp_p_6/out_left.n1 comp_p_6/out_left.t2 145.612
R3729 comp_p_6/out_left.n2 comp_p_6/out_left.t0 143.417
R3730 comp_p_6/out_left.n0 comp_p_6/out_left.t1 29.4286
R3731 comp_p_6/out_left comp_p_6/out_left.n3 11.6041
R3732 comp_p_6/out_left.n3 comp_p_6/out_left.n2 4.33076
R3733 comp_p_6/out_left.n1 comp_p_6/out_left.n0 2.12634
R3734 comp_p_6/out_left.n2 comp_p_6/out_left.n1 2.04428
R3735 comp_p_6/out_left.n3 comp_p_6/out_left.n0 0.00290385
R3736 d6.n0 d6.t1 556.78
R3737 d6.t1 d6 547.24
R3738 d6 d6.t0 372.113
R3739 d6.n1 d6 11.4942
R3740 d6.n0 d6 9.54008
R3741 d6.n3 d6 7.39314
R3742 d6.n2 d6.n1 3.43599
R3743 d6.n1 d6 1.33473
R3744 d6 d6.n3 0.714431
R3745 d6 d6.n0 0.266125
R3746 d6 d6 0.063
R3747 d6.n3 d6 0.0550806
R3748 d6.n3 d6.n2 0.00313551
R3749 d6.n2 d6 0.00313551
R3750 dout0 dout0 5.30089
R3751 dout0 dout0 2.61734
R3752 dout1 dout1 5.30089
R3753 dout1 dout1 2.61734
R3754 dout2 dout2 5.30089
R3755 dout2 dout2 2.61734
C0 vdd comp_p_0/out_left 0.01217f
C1 comp_p_6/latch_left d4 0.06068f
C2 comp_p_2/vinn comp_p_2/tail 0
C3 comp_p_6/vbias_p comp_p_2/latch_right 0.40389f
C4 vbias_generation_0/bias_n comp_p_6/vbias_p 0
C5 vbias_generation_0/XR_bias_4/R1 comp_p_6/vinn 0.51064f
C6 comp_p_4/tail comp_p_5/vinn 0.10856f
C7 vdd comp_p_1/latch_left 2.04615f
C8 comp_p_1/vinn comp_p_0/vinn 0.94729f
C9 d4 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C10 tmux_7therm_to_3bin_0/buffer_5/out d4 0.01353f
C11 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d6 0
C12 vin comp_p_2/latch_right 0.21614f
C13 d5 d0 0.04762f
C14 d2 tmux_7therm_to_3bin_0/R1/R1 0.00763f
C15 vbias_generation_0/bias_n vin 0.0214f
C16 tmux_7therm_to_3bin_0/buffer_4/out vdd 0.00846f
C17 d5 comp_p_1/out_left 0
C18 comp_p_6/vbias_p comp_p_4/vinn 0.12306f
C19 vbias_generation_0/XR_bias_2/R2 comp_p_6/vinn 0.00358f
C20 d2 tmux_7therm_to_3bin_0/buffer_1/out 0
C21 d5 comp_p_3/out_left 0.02324f
C22 comp_p_6/tail d4 0.00252f
C23 d2 comp_p_1/latch_right 0.00123f
C24 vin d6 0.01178f
C25 comp_p_4/latch_left comp_p_5/vinn 0.16266f
C26 d5 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C27 comp_p_5/tail vdd 0.35567f
C28 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d4 0.00318f
C29 vbias_generation_0/XR_bias_4/R1 comp_p_4/latch_right 0
C30 vin comp_p_4/vinn 0.52728f
C31 d4 comp_p_6/vbias_p 0.37293f
C32 comp_p_0/latch_right d1 0
C33 comp_p_6/out_left vbias_generation_0/bias_n 0.00925f
C34 d5 comp_p_3/vinn 0
C35 d5 d3 0.16529f
C36 tmux_7therm_to_3bin_0/buffer_0/out vdd 0
C37 d5 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.00186f
C38 d4 vin 0.72855f
C39 d2 tmux_7therm_to_3bin_0/buffer_2/out 0
C40 comp_p_2/vinn comp_p_0/vinn 0.02754f
C41 d2 vdd 1.1602f
C42 comp_p_4/out_left comp_p_4/vinn 0.02516f
C43 d5 comp_p_1/latch_left 0
C44 comp_p_6/latch_left vin 0.00266f
C45 vdd comp_p_5/latch_right 1.9557f
C46 comp_p_6/out_left d4 0.27385f
C47 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vdd 0
C48 vdd comp_p_2/tail 0.00168f
C49 d5 tmux_7therm_to_3bin_0/buffer_4/out 0
C50 comp_p_5/out_left comp_p_4/tail 0
C51 d1 comp_p_2/latch_right 0.01472f
C52 vdd tmux_7therm_to_3bin_0/tmux_2to1_3/A 0.00153f
C53 comp_p_0/latch_right comp_p_1/out_left 0
C54 vdd comp_p_4/tail 0.00166f
C55 vbias_generation_0/bias_n comp_p_6/vinn 0.43753f
C56 comp_p_6/tail vin 0
C57 comp_p_2/out_left comp_p_3/vinn 0.01462f
C58 d1 d6 0.09f
C59 vdd tmux_7therm_to_3bin_0/buffer_8/in 0
C60 vin comp_p_6/vbias_p 1.44761f
C61 tmux_7therm_to_3bin_0/buffer_0/out d5 0
C62 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d6 0.00531f
C63 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin vdd 0.00196f
C64 comp_p_2/out_left comp_p_0/out_left 0.09264f
C65 d2 d5 0.04508f
C66 vdd comp_p_1/tail 0.35563f
C67 comp_p_0/vinn comp_p_2/latch_left 0
C68 d4 d1 0.33457f
C69 vdd comp_p_4/latch_left 0
C70 comp_p_6/out_left comp_p_6/vbias_p -0.05282f
C71 d2 comp_p_3/tail 0.00272f
C72 vbias_generation_0/bias_n comp_p_4/latch_right 0
C73 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d4 0.00248f
C74 vdd comp_p_0/vinn 0.01961f
C75 d4 comp_p_6/vinn 0.06841f
C76 comp_p_6/vbias_p comp_p_4/out_left 0.69034f
C77 comp_p_0/latch_right comp_p_1/latch_left 0.02598f
C78 comp_p_6/out_left vin 0.06197f
C79 comp_p_6/latch_left comp_p_6/vinn 0.00473f
C80 comp_p_4/latch_right comp_p_4/vinn 0.00144f
C81 comp_p_1/latch_right comp_p_1/vinn 0.00799f
C82 comp_p_2/latch_right comp_p_3/out_left 0
C83 vin comp_p_4/out_left 0.0859f
C84 dout0 dout1 -0
C85 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d1 0.00173f
C86 d0 d6 0.09283f
C87 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin tmux_7therm_to_3bin_0/R1/R1 0
C88 comp_p_1/out_left d6 0
C89 comp_p_0/tail comp_p_1/vinn 0.10698f
C90 d4 comp_p_4/latch_right 0
C91 d6 comp_p_3/out_left 0
C92 tmux_7therm_to_3bin_0/R1/m1_n100_n100# d3 0
C93 comp_p_1/vinn comp_p_2/latch_left 0.01672f
C94 comp_p_3/vinn comp_p_2/latch_right 0.17593f
C95 d6 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C96 d5 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C97 vdd comp_p_1/vinn 1.45687f
C98 d4 d0 0.03391f
C99 vdd comp_p_6/latch_right 1.95582f
C100 d5 comp_p_1/tail 0
C101 comp_p_6/vbias_p d1 0.37529f
C102 d4 comp_p_1/out_left 0
C103 vbias_generation_0/XR_bias_3/R2 comp_p_6/tail 0
C104 d6 comp_p_3/vinn 0
C105 d4 comp_p_3/out_left 0
C106 d3 d6 0.07956f
C107 comp_p_6/vbias_p comp_p_6/vinn 0.31983f
C108 d2 comp_p_0/latch_right 0.01472f
C109 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d6 0
C110 comp_p_5/out_left comp_p_5/vinn 0.19629f
C111 comp_p_3/vinn comp_p_4/vinn 0
C112 d4 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C113 vin d1 0.63586f
C114 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin vdd 0
C115 vref vin 0.00582f
C116 comp_p_1/latch_right comp_p_3/latch_right 0.00925f
C117 vbias_generation_0/XR_bias_3/R2 vin 0.08368f
C118 vin comp_p_6/vinn 1.01745f
C119 d4 comp_p_3/vinn 0
C120 comp_p_3/latch_left vdd 2.04611f
C121 d6 comp_p_1/latch_left 0
C122 vdd comp_p_5/vinn 1.45079f
C123 d4 d3 2.88908f
C124 d4 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.00384f
C125 comp_p_2/vinn comp_p_2/latch_left 0
C126 vbias_generation_0/XR_bias_4/R1 comp_p_4/latch_left 0
C127 tmux_7therm_to_3bin_0/buffer_4/out d6 0
C128 comp_p_6/vbias_p comp_p_4/latch_right 0.40389f
C129 vdd comp_p_2/vinn 0.04727f
C130 vbias_generation_0/XR_bias_3/R2 comp_p_6/out_left 0.00563f
C131 comp_p_6/out_left comp_p_6/vinn 0.14972f
C132 vdd comp_p_3/latch_right 1.95698f
C133 d4 comp_p_1/latch_left 0
C134 tmux_7therm_to_3bin_0/R1/R1 tmux_7therm_to_3bin_0/buffer_1/out 0
C135 d0 comp_p_6/vbias_p 0.00465f
C136 comp_p_6/vinn comp_p_4/out_left 0.04948f
C137 comp_p_5/tail d6 0
C138 vin comp_p_4/latch_right 0.21628f
C139 d5 comp_p_1/vinn 0
C140 comp_p_6/vbias_p comp_p_1/out_left -0.065f
C141 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d3 0
C142 d4 tmux_7therm_to_3bin_0/buffer_4/out 0
C143 tmux_7therm_to_3bin_0/R1/R2 d3 0
C144 comp_p_5/latch_left comp_p_5/vinn 0.00674f
C145 d2 comp_p_2/latch_right 0.00137f
C146 comp_p_6/vbias_p comp_p_3/out_left -0.06014f
C147 tmux_7therm_to_3bin_0/buffer_0/out d6 0
C148 comp_p_2/out_left comp_p_0/vinn 0.0271f
C149 vin comp_p_1/out_left 0.07139f
C150 comp_p_5/tail d4 0.00264f
C151 d2 d6 0.05303f
C152 vin comp_p_3/out_left 0.05071f
C153 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d5 0
C154 tmux_7therm_to_3bin_0/R1/R1 vdd 0.00399f
C155 vdd tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G 0.00166f
C156 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d3 0
C157 comp_p_6/vbias_p comp_p_3/vinn 0.38072f
C158 d3 comp_p_6/vbias_p 0
C159 comp_p_0/latch_right comp_p_0/vinn 0.00236f
C160 comp_p_3/latch_left d5 0
C161 comp_p_5/latch_right d6 0
C162 tmux_7therm_to_3bin_0/buffer_0/out d4 0
C163 comp_p_6/vbias_p comp_p_0/out_left 0.68459f
C164 comp_p_1/latch_right vdd 1.96641f
C165 vin comp_p_3/vinn 0.65736f
C166 d2 d4 0.04942f
C167 vin d3 0.00158f
C168 vref comp_p_6/vinn 0.00148f
C169 comp_p_5/out_left vdd 1.8042f
C170 vbias_generation_0/XR_bias_3/R2 comp_p_6/vinn 0.06411f
C171 comp_p_0/tail vdd 0.00166f
C172 d5 comp_p_3/latch_right 0.00185f
C173 vin comp_p_0/out_left 0.0787f
C174 d4 comp_p_5/latch_right 0.06539f
C175 vdd comp_p_2/latch_left 0
C176 comp_p_0/latch_left comp_p_0/vinn 0.02494f
C177 comp_p_2/out_left comp_p_1/vinn 0.00265f
C178 d2 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0.00483f
C179 comp_p_0/latch_right comp_p_1/vinn 0.1958f
C180 vbias_generation_0/bias_n comp_p_4/latch_left 0
C181 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d6 0
C182 comp_p_6/vinn comp_p_4/latch_right 0.00583f
C183 d4 comp_p_4/tail -0.00224f
C184 comp_p_1/tail d6 0
C185 d0 d1 1.12322f
C186 comp_p_1/out_left d1 0.67001f
C187 comp_p_5/tail vin 0.00233f
C188 comp_p_4/latch_left comp_p_4/vinn 0.00288f
C189 comp_p_5/latch_left vdd 2.0461f
C190 d2 comp_p_6/vbias_p 0.37534f
C191 comp_p_0/latch_left comp_p_1/vinn 0.15776f
C192 d4 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C193 comp_p_1/latch_right d5 0.0019f
C194 comp_p_2/out_left comp_p_2/vinn 0.0232f
C195 d4 comp_p_1/tail 0
C196 comp_p_5/out_left d5 0
C197 d2 vin 0.72189f
C198 d1 comp_p_3/vinn 0
C199 d3 d1 0.11517f
C200 comp_p_6/vbias_p comp_p_2/tail 0.31443f
C201 d5 vdd 2.33637f
C202 comp_p_1/vinn comp_p_2/latch_right 0.00771f
C203 vbias_generation_0/bias_n comp_p_6/latch_right 0
C204 vin comp_p_2/tail 0.0104f
C205 d1 comp_p_1/latch_left 0.09502f
C206 comp_p_3/tail vdd 0.35691f
C207 comp_p_4/tail comp_p_6/vbias_p 0.31443f
C208 d6 comp_p_1/vinn 0
C209 d0 comp_p_1/out_left -0
C210 vin comp_p_4/tail 0.01181f
C211 comp_p_3/latch_left comp_p_2/latch_right 0.02598f
C212 d4 comp_p_1/vinn 0
C213 d4 comp_p_6/latch_right 0.06065f
C214 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d6 0
C215 comp_p_6/vbias_p comp_p_4/latch_left 0.37827f
C216 d0 d3 0.03225f
C217 d6 comp_p_5/vinn 0.00513f
C218 comp_p_2/vinn comp_p_2/latch_right 0
C219 comp_p_3/latch_left d6 0
C220 d3 comp_p_1/out_left 0
C221 comp_p_6/vbias_p comp_p_0/vinn 0.12305f
C222 comp_p_3/vinn comp_p_3/out_left 0.20126f
C223 vin comp_p_1/tail 0.00233f
C224 comp_p_5/vinn comp_p_4/vinn 0.32186f
C225 tmux_7therm_to_3bin_0/buffer_0/out d1 0
C226 vin comp_p_4/latch_left 0.00664f
C227 comp_p_2/out_left vdd 0.02487f
C228 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d4 0
C229 d2 d1 3.44306f
C230 d3 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0.00238f
C231 vin comp_p_0/vinn 0.81463f
C232 d6 comp_p_3/latch_right 0.00265f
C233 comp_p_3/latch_left d4 0
C234 d4 comp_p_5/vinn 0.25734f
C235 comp_p_0/latch_right vdd 0.00588f
C236 comp_p_3/tail d5 0
C237 d3 comp_p_3/vinn 0.0076f
C238 d4 comp_p_3/latch_right 0.00133f
C239 comp_p_0/latch_left comp_p_2/latch_left 0.01494f
C240 comp_p_6/vbias_p comp_p_1/vinn 0.38594f
C241 d3 comp_p_1/latch_left 0
C242 comp_p_0/latch_left vdd 0
C243 tmux_7therm_to_3bin_0/buffer_6/out d6 0
C244 vin comp_p_1/vinn 0.97735f
C245 tmux_7therm_to_3bin_0/buffer_0/out d0 0
C246 d2 d0 0.03281f
C247 comp_p_1/latch_right d6 0.00271f
C248 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d1 0.00131f
C249 d2 comp_p_1/out_left 0
C250 tmux_7therm_to_3bin_0/R1/R1 d4 0
C251 d2 comp_p_3/out_left 0.67197f
C252 d4 tmux_7therm_to_3bin_0/buffer_6/out 0.013f
C253 comp_p_5/out_left d6 0
C254 comp_p_6/vbias_p comp_p_5/vinn 0.407f
C255 vdd comp_p_2/latch_right 0.00592f
C256 d1 comp_p_1/tail 0.00457f
C257 vbias_generation_0/bias_n vdd 0.0189f
C258 d4 tmux_7therm_to_3bin_0/buffer_1/out 0
C259 comp_p_5/out_left comp_p_4/vinn 0
C260 comp_p_1/latch_right d4 0
C261 d1 comp_p_0/vinn -0
C262 comp_p_4/latch_left comp_p_6/vinn 0.00606f
C263 vin comp_p_5/vinn 0.66275f
C264 tmux_7therm_to_3bin_0/buffer_0/out d3 0
C265 comp_p_6/vbias_p comp_p_2/vinn 0.12413f
C266 vdd d6 5.14819f
C267 d2 comp_p_3/vinn 0.24742f
C268 comp_p_5/out_left d4 0.61081f
C269 d2 d3 2.50136f
C270 vdd comp_p_4/vinn 0.03662f
C271 comp_p_2/tail comp_p_3/out_left 0
C272 d0 tmux_7therm_to_3bin_0/tmux_2to1_3/A 0
C273 vin comp_p_2/vinn 0.52215f
C274 tmux_7therm_to_3bin_0/buffer_2/out d4 0
C275 d4 vdd 1.46527f
C276 d2 comp_p_1/latch_left 0
C277 m3_n3070_n10912# vin 0.06232f
C278 comp_p_2/tail comp_p_3/vinn 0.14685f
C279 comp_p_5/vinn comp_p_4/out_left 0.01843f
C280 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d0 0.00746f
C281 comp_p_5/latch_left d6 0.00183f
C282 comp_p_6/latch_left vdd 2.04625f
C283 d1 comp_p_1/vinn 0.26331f
C284 comp_p_6/latch_right comp_p_6/vinn 0.00296f
C285 comp_p_1/out_left comp_p_0/vinn 0
C286 comp_p_5/latch_left d4 0.06545f
C287 d5 d6 4.44886f
C288 comp_p_5/out_left comp_p_6/vbias_p -0.0642f
C289 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d3 0
C290 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d1 0.00482f
C291 comp_p_0/tail comp_p_6/vbias_p 0.31443f
C292 comp_p_6/vbias_p comp_p_2/latch_left 0.37827f
C293 d2 tmux_7therm_to_3bin_0/buffer_0/out 0
C294 comp_p_6/tail vdd 0.35623f
C295 d3 comp_p_1/tail 0
C296 comp_p_6/latch_left comp_p_5/latch_left 0.00925f
C297 comp_p_3/latch_left d1 0
C298 comp_p_3/tail d6 0
C299 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vdd 0.00104f
C300 comp_p_5/out_left vin 0.06043f
C301 comp_p_0/latch_left comp_p_2/out_left 0.01472f
C302 vdd comp_p_6/vbias_p 12.48384f
C303 comp_p_0/tail vin 0.01181f
C304 comp_p_3/vinn comp_p_0/vinn 0.53686f
C305 comp_p_6/vinn comp_p_5/vinn 0.03037f
C306 d4 d5 4.51321f
C307 vin comp_p_2/latch_left 0.00664f
C308 comp_p_0/out_left comp_p_0/vinn 0.02276f
C309 d1 comp_p_3/latch_right 0
C310 vin vdd 10.39915f
C311 comp_p_3/tail d4 0
C312 d2 comp_p_2/tail -0.00224f
C313 comp_p_1/out_left comp_p_1/vinn 0.19389f
C314 vref m3_n3070_n10912# 0.5517f
C315 m3_n3070_n10912# comp_p_6/vinn 0.08555f
C316 comp_p_6/out_left vdd 1.84652f
C317 d5 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C318 comp_p_5/vinn comp_p_4/latch_right 0.20935f
C319 tmux_7therm_to_3bin_0/buffer_5/out d5 0
C320 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d0 0
C321 comp_p_0/latch_right comp_p_2/latch_right 0.01494f
C322 vdd comp_p_4/out_left 0.02489f
C323 comp_p_1/vinn comp_p_3/vinn 0.03321f
C324 d3 comp_p_1/vinn 0
C325 tmux_7therm_to_3bin_0/R1/R1 d1 0.00785f
C326 d2 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C327 d1 tmux_7therm_to_3bin_0/buffer_1/out 0.01311f
C328 comp_p_1/vinn comp_p_0/out_left 0.04644f
C329 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d5 0
C330 d5 comp_p_6/vbias_p 0
C331 d2 comp_p_1/tail 0
C332 comp_p_1/latch_right d1 0.09536f
C333 comp_p_1/vinn comp_p_1/latch_left 0.0067f
C334 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d3 0
C335 comp_p_2/vinn comp_p_3/out_left 0
C336 comp_p_0/tail d1 -0.00224f
C337 d5 vin 0.0056f
C338 comp_p_5/vinn comp_p_3/vinn 0.0226f
C339 comp_p_3/latch_left comp_p_3/vinn 0.00666f
C340 comp_p_3/latch_left d3 0
C341 tmux_7therm_to_3bin_0/buffer_2/out d1 0.00551f
C342 comp_p_3/tail vin 0.00233f
C343 vdd d1 1.15842f
C344 comp_p_2/vinn comp_p_3/vinn 0.31389f
C345 vbias_generation_0/XR_bias_4/R1 comp_p_6/vbias_p 0.02724f
C346 vref vdd 0
C347 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin vdd 0.00122f
C348 vbias_generation_0/XR_bias_3/R2 vdd 0.08059f
C349 vdd comp_p_6/vinn 1.11418f
C350 comp_p_3/vinn comp_p_3/latch_right 0.00805f
C351 comp_p_3/latch_left comp_p_1/latch_left 0.00925f
C352 d3 comp_p_3/latch_right 0.0057f
C353 tmux_7therm_to_3bin_0/R1/R1 d0 0.00538f
C354 d0 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G 0
C355 vbias_generation_0/XR_bias_4/R1 vin 0.00472f
C356 vbias_generation_0/XR_bias_2/R2 comp_p_6/vbias_p 0.02749f
C357 comp_p_5/out_left comp_p_4/latch_right 0
C358 d2 comp_p_1/vinn 0.00152f
C359 comp_p_2/out_left comp_p_6/vbias_p 0.68901f
C360 vbias_generation_0/XR_bias_2/R2 vin 0.50675f
C361 vdd comp_p_4/latch_right 0.00589f
C362 comp_p_5/latch_right comp_p_6/latch_right 0.00925f
C363 comp_p_0/tail comp_p_1/out_left 0
C364 d4 vbias_generation_0/bias_n 0.00802f
C365 tmux_7therm_to_3bin_0/R1/R1 d3 0
C366 comp_p_2/out_left vin 0.0842f
C367 comp_p_5/out_left comp_p_3/out_left 0.01584f
C368 comp_p_0/latch_right comp_p_6/vbias_p 0.40389f
C369 vbias_generation_0/XR_bias_4/R1 comp_p_4/out_left 0
C370 d3 tmux_7therm_to_3bin_0/buffer_1/out 0
C371 d2 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0.00171f
C372 d0 vdd 2.71992f
C373 d4 d6 0.79887f
C374 vdd comp_p_1/out_left 1.79183f
C375 comp_p_1/latch_right d3 0.00104f
C376 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vdd 0.00166f
C377 comp_p_6/latch_left vbias_generation_0/bias_n 0.01259f
C378 d2 comp_p_3/latch_left 0.09614f
C379 comp_p_0/latch_right vin 0.21598f
C380 d5 d1 0.26099f
C381 d4 comp_p_4/vinn -0
C382 vdd comp_p_3/out_left 1.79594f
C383 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d5 0
C384 comp_p_5/out_left d3 0.02309f
C385 vdd tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C386 comp_p_0/latch_left comp_p_6/vbias_p 0.37827f
C387 comp_p_3/vinn comp_p_2/latch_left 0.15548f
C388 comp_p_5/latch_right comp_p_5/vinn 0.00802f
C389 comp_p_5/latch_left comp_p_4/latch_right 0.02598f
C390 comp_p_2/out_left comp_p_4/out_left 0.01584f
C391 d2 comp_p_3/latch_right 0.09517f
C392 vdd comp_p_3/vinn 1.48772f
C393 tmux_7therm_to_3bin_0/buffer_2/out d3 0
C394 comp_p_0/out_left comp_p_2/latch_left 0.01472f
C395 vdd d3 2.3721f
C396 comp_p_0/latch_left vin 0.00334f
C397 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin vdd 0.00104f
C398 vdd tmux_7therm_to_3bin_0/buffer_7/in 0.0027f
C399 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d6 0
C400 m3_n3070_n10912# vss 0.95701f $ **FLOATING
C401 d6.t1 vss 0.09646f
C402 d6.t0 vss 0.09152f
C403 d6.n0 vss 0.27307f
C404 d6.n1 vss 2.87854f
C405 d6.n2 vss 0.46328f
C406 d6.n3 vss 28.1493f
C407 comp_p_6/out_left.t1 vss 0.35725f
C408 comp_p_6/out_left.n0 vss 0.35824f
C409 comp_p_6/out_left.t2 vss 0.95164f
C410 comp_p_6/out_left.n1 vss 1.72525f
C411 comp_p_6/out_left.t0 vss 0.94389f
C412 comp_p_6/out_left.n2 vss 0.3128f
C413 comp_p_6/out_left.n3 vss 1.23781f
C414 comp_p_6/latch_left.t0 vss 1.25281f
C415 comp_p_6/latch_left.t3 vss 1.57061f
C416 comp_p_6/latch_left.t2 vss 1.45859f
C417 comp_p_6/latch_left.n0 vss 2.77309f
C418 comp_p_6/latch_left.n1 vss 1.77973f
C419 comp_p_6/latch_left.t1 vss 0.37457f
C420 comp_p_6/latch_left.n2 vss 1.60078f
C421 d5.t0 vss 0.55064f
C422 d5.t1 vss 0.58031f
C423 d5.n0 vss 1.64287f
C424 d5.n1 vss 4.12658f
C425 comp_p_5/latch_left.t0 vss 1.25281f
C426 comp_p_5/latch_left.t3 vss 1.57061f
C427 comp_p_5/latch_left.t2 vss 1.45859f
C428 comp_p_5/latch_left.n0 vss 2.77309f
C429 comp_p_5/latch_left.n1 vss 1.77973f
C430 comp_p_5/latch_left.t1 vss 0.37457f
C431 comp_p_5/latch_left.n2 vss 1.60078f
C432 d4.t1 vss 0.06875f
C433 d4.t0 vss 0.06524f
C434 d4.n0 vss 0.19465f
C435 d4.n1 vss 4.22355f
C436 d4.n2 vss 6.74001f
C437 comp_p_4/out_left.t1 vss 0.26539f
C438 comp_p_4/out_left.n0 vss 0.26612f
C439 comp_p_4/out_left.t2 vss 0.70693f
C440 comp_p_4/out_left.n1 vss 1.28162f
C441 comp_p_4/out_left.t0 vss 0.70117f
C442 comp_p_4/out_left.n2 vss 0.23237f
C443 comp_p_4/out_left.n3 vss 0.91952f
C444 comp_p_4/latch_left.t0 vss 1.01079f
C445 comp_p_4/latch_left.t3 vss 1.2672f
C446 comp_p_4/latch_left.t2 vss 1.17681f
C447 comp_p_4/latch_left.n0 vss 2.23738f
C448 comp_p_4/latch_left.n1 vss 1.43592f
C449 comp_p_4/latch_left.t1 vss 0.30221f
C450 comp_p_4/latch_left.n2 vss 1.29154f
C451 d3.t0 vss 0.10693f
C452 d3.t1 vss 0.11269f
C453 d3.n0 vss 0.31904f
C454 d3.n1 vss 2.47445f
C455 d3.n2 vss 0.38144f
C456 d3.n3 vss 7.05226f
C457 comp_p_3/out_left.t1 vss 0.35725f
C458 comp_p_3/out_left.n0 vss 0.35824f
C459 comp_p_3/out_left.t2 vss 0.95164f
C460 comp_p_3/out_left.n1 vss 1.72525f
C461 comp_p_3/out_left.t0 vss 0.94389f
C462 comp_p_3/out_left.n2 vss 0.3128f
C463 comp_p_3/out_left.n3 vss 1.23781f
C464 comp_p_3/latch_right.t1 vss 0.4606f
C465 comp_p_3/latch_right.n0 vss 0.90852f
C466 comp_p_3/latch_right.t3 vss 1.93136f
C467 comp_p_3/latch_right.t2 vss 1.7936f
C468 comp_p_3/latch_right.n1 vss 3.06813f
C469 comp_p_3/latch_right.t0 vss 1.53795f
C470 comp_p_3/latch_right.n2 vss 0.44996f
C471 comp_p_3/latch_right.n3 vss 2.026f
C472 comp_p_3/latch_right.n4 vss 0.28331f
C473 comp_p_3/latch_left.t0 vss 1.25281f
C474 comp_p_3/latch_left.t3 vss 1.57061f
C475 comp_p_3/latch_left.t2 vss 1.45859f
C476 comp_p_3/latch_left.n0 vss 2.77309f
C477 comp_p_3/latch_left.n1 vss 1.77973f
C478 comp_p_3/latch_left.t1 vss 0.37457f
C479 comp_p_3/latch_left.n2 vss 1.60078f
C480 d2.t1 vss 0.08206f
C481 d2.t0 vss 0.07786f
C482 d2.n0 vss 0.23064f
C483 d2.n1 vss 0.05046f
C484 d2.n2 vss 3.22714f
C485 d2.n3 vss 0.16699f
C486 d2.n4 vss 6.27226f
C487 comp_p_2/latch_left.t0 vss 1.01079f
C488 comp_p_2/latch_left.t3 vss 1.2672f
C489 comp_p_2/latch_left.t2 vss 1.17681f
C490 comp_p_2/latch_left.n0 vss 2.23738f
C491 comp_p_2/latch_left.n1 vss 1.43592f
C492 comp_p_2/latch_left.t1 vss 0.30221f
C493 comp_p_2/latch_left.n2 vss 1.29154f
C494 d1.t0 vss 0.05868f
C495 d1.t1 vss 0.06184f
C496 d1.n0 vss 0.17507f
C497 d1.n1 vss 2.81604f
C498 d1.n2 vss 1.53469f
C499 comp_p_0/out_left.t1 vss 0.26539f
C500 comp_p_0/out_left.n0 vss 0.26612f
C501 comp_p_0/out_left.t2 vss 0.70693f
C502 comp_p_0/out_left.n1 vss 1.28162f
C503 comp_p_0/out_left.t0 vss 0.70117f
C504 comp_p_0/out_left.n2 vss 0.23237f
C505 comp_p_0/out_left.n3 vss 0.91952f
C506 vin.t4 vss 0.59319f
C507 vin.t5 vss 0.5928f
C508 vin.n0 vss 0.79649f
C509 vin.n1 vss 0.62357f
C510 vin.t6 vss 0.44086f
C511 vin.n2 vss 0.7172f
C512 vin.t7 vss 0.4403f
C513 vin.n3 vss 0.70513f
C514 vin.n4 vss 0.3342f
C515 vin.t8 vss 0.59319f
C516 vin.t9 vss 0.5928f
C517 vin.n5 vss 0.79649f
C518 vin.n6 vss 0.62357f
C519 vin.t10 vss 0.44086f
C520 vin.n7 vss 0.7172f
C521 vin.t11 vss 0.4403f
C522 vin.n8 vss 0.70513f
C523 vin.n9 vss 0.3342f
C524 vin.n10 vss 4.90773f
C525 vin.t16 vss 0.59319f
C526 vin.t17 vss 0.5928f
C527 vin.n11 vss 0.79649f
C528 vin.n12 vss 0.62357f
C529 vin.t18 vss 0.44086f
C530 vin.n13 vss 0.7172f
C531 vin.t19 vss 0.4403f
C532 vin.n14 vss 0.70513f
C533 vin.n15 vss 0.3342f
C534 vin.n16 vss 2.83617f
C535 vin.n17 vss 1.64566f
C536 vin.t24 vss 0.59319f
C537 vin.t25 vss 0.5928f
C538 vin.n18 vss 0.79649f
C539 vin.n19 vss 0.62357f
C540 vin.t26 vss 0.44086f
C541 vin.n20 vss 0.7172f
C542 vin.t27 vss 0.4403f
C543 vin.n21 vss 0.70513f
C544 vin.n22 vss 0.3342f
C545 vin.t0 vss 0.59319f
C546 vin.t1 vss 0.5928f
C547 vin.n23 vss 0.79649f
C548 vin.n24 vss 0.62357f
C549 vin.t2 vss 0.44086f
C550 vin.n25 vss 0.7172f
C551 vin.t3 vss 0.4403f
C552 vin.n26 vss 0.70513f
C553 vin.n27 vss 0.32342f
C554 vin.n28 vss 1.51786f
C555 vin.t12 vss 0.59319f
C556 vin.t13 vss 0.5928f
C557 vin.n29 vss 0.79649f
C558 vin.n30 vss 0.62357f
C559 vin.t14 vss 0.44086f
C560 vin.n31 vss 0.7172f
C561 vin.t15 vss 0.4403f
C562 vin.n32 vss 0.70513f
C563 vin.n33 vss 0.33241f
C564 vin.n34 vss 0.34098f
C565 vin.n35 vss 5.06577f
C566 vin.t20 vss 0.59319f
C567 vin.t21 vss 0.5928f
C568 vin.n36 vss 0.79649f
C569 vin.n37 vss 0.62357f
C570 vin.t22 vss 0.44086f
C571 vin.n38 vss 0.7172f
C572 vin.t23 vss 0.4403f
C573 vin.n39 vss 0.70513f
C574 vin.n40 vss 0.3265f
C575 vin.n41 vss 0.44248f
C576 vin.n42 vss 3.93947f
C577 vin.n43 vss 3.62493f
C578 vin.n44 vss 1.93496f
C579 vin.n45 vss 1.86174f
C580 d0.t1 vss 0.07597f
C581 d0.t0 vss 0.07208f
C582 d0.n0 vss 0.21301f
C583 d0.n1 vss 0.04873f
C584 d0.n2 vss 1.26804f
C585 d0.n3 vss 0.90329f
C586 comp_p_1/latch_left.t0 vss 1.25281f
C587 comp_p_1/latch_left.t3 vss 1.57061f
C588 comp_p_1/latch_left.t2 vss 1.45859f
C589 comp_p_1/latch_left.n0 vss 2.77309f
C590 comp_p_1/latch_left.n1 vss 1.77973f
C591 comp_p_1/latch_left.t1 vss 0.37457f
C592 comp_p_1/latch_left.n2 vss 1.60078f
C593 vdd.n0 vss 2.61314f
C594 vdd.n1 vss 0.35701f
C595 vdd.n2 vss 0.25978f
C596 vdd.n3 vss 0.3522f
C597 vdd.n4 vss 0.06614f
C598 vdd.n5 vss 0.41889f
C599 vdd.n6 vss 0.5445f
C600 vdd.n7 vss 0.02158f
C601 vdd.n8 vss 0.14159f
C602 vdd.n9 vss 0.03904f
C603 vdd.n10 vss 0.02097f
C604 vdd.n11 vss 1.37952f
C605 vdd.n12 vss 0.05232f
C606 vdd.n13 vss 0.05047f
C607 vdd.n14 vss 0.96343f
C608 vdd.n15 vss 0.05028f
C609 vdd.n16 vss 1.20937f
C610 vdd.n17 vss 0.35256f
C611 vdd.n18 vss 0.13091f
C612 vdd.n19 vss 1.10027f
C613 vdd.n20 vss 0.75668f
C614 vdd.n21 vss 0.22818f
C615 vdd.n22 vss 0.79714f
C616 vdd.n23 vss 0.29863f
C617 vdd.n24 vss 0.04637f
C618 vdd.n25 vss 0.05028f
C619 vdd.n26 vss 0.06016f
C620 vdd.n27 vss 0.04638f
C621 vdd.n28 vss 1.10725f
C622 vdd.n29 vss 1.55964f
C623 vdd.n30 vss 0.44293f
C624 vdd.n31 vss 0.11722f
C625 vdd.n32 vss 0.16179f
C626 vdd.n33 vss 0.03916f
C627 vdd.n34 vss 0.03615f
C628 vdd.n35 vss 0.27022f
C629 vdd.n36 vss 0.81131f
C630 vdd.n37 vss 0.25716f
C631 vdd.n38 vss 1.575f
C632 vdd.n39 vss 0.05047f
C633 vdd.n40 vss 0.05047f
C634 vdd.n41 vss 0.83064f
C635 vdd.n42 vss 0.04638f
C636 vdd.n43 vss 0.14124f
C637 vdd.n44 vss 0.05028f
C638 vdd.n45 vss 0.05028f
C639 vdd.n46 vss 1.34881f
C640 vdd.n47 vss 1.58198f
C641 vdd.n48 vss 0.03904f
C642 vdd.n49 vss 0.03904f
C643 vdd.n50 vss 0.02158f
C644 vdd.n51 vss -0.10005f
C645 vdd.n52 vss 0.05057f
C646 vdd.n53 vss 0.0514f
C647 vdd.n54 vss 0.02369f
C648 vdd.n55 vss 1.21001f
C649 vdd.n56 vss 1.10725f
C650 vdd.n57 vss 0.05045f
C651 vdd.n58 vss 0.13743f
C652 vdd.n59 vss 0.03916f
C653 vdd.n60 vss 1.6455f
C654 vdd.n61 vss 0.04413f
C655 vdd.n62 vss 0.27022f
C656 vdd.n63 vss 0.44293f
C657 vdd.n64 vss 0.81131f
C658 vdd.n65 vss 0.25716f
C659 vdd.n66 vss 0.03615f
C660 vdd.n67 vss 0.03916f
C661 vdd.n68 vss 1.55964f
C662 vdd.n69 vss 0.30997f
C663 vdd.n70 vss 0.05045f
C664 vdd.n71 vss 0.13183f
C665 vdd.n72 vss 0.13091f
C666 vdd.n73 vss 0.05057f
C667 vdd.n74 vss 0.24854f
C668 vdd.n75 vss 1.11563f
C669 vdd.n76 vss 0.0514f
C670 vdd.n77 vss 0.45695f
C671 vdd.n78 vss 0.00715f
C672 vdd.n79 vss 0.14251f
C673 vdd.n80 vss 0.03916f
C674 vdd.n81 vss 4.65538f
C675 vdd.n82 vss 0.1416f
C676 vdd.n83 vss 0.00288f
C677 vdd.n84 vss 0.01263f
C678 vdd.n85 vss 0.01873f
C679 vdd.n86 vss 0.01203f
C680 vdd.n87 vss 0.01873f
C681 vdd.n88 vss 0.14091f
C682 vdd.n89 vss 0.01263f
C683 vdd.n90 vss 0.01203f
C684 vdd.n91 vss 0.01203f
C685 vdd.n92 vss 0.01203f
C686 vdd.n93 vss 0.14091f
C687 vdd.n94 vss 0.01245f
C688 vdd.n95 vss 0.01245f
C689 vdd.n96 vss 0.14091f
C690 vdd.n97 vss 0.01919f
C691 vdd.n98 vss 0.01919f
C692 vdd.n99 vss 0.0067f
C693 vdd.n100 vss 0.00961f
C694 vdd.n101 vss 0.15437f
C695 vdd.n102 vss 0.01919f
C696 vdd.n103 vss 0.01919f
C697 vdd.n104 vss 0.08965f
C698 vdd.n105 vss 0.05327f
C699 vdd.n106 vss 0.17275f
C700 vdd.n107 vss 0.00944f
C701 vdd.n108 vss 0.00961f
C702 vdd.n110 vss 0.12299f
C703 vdd.n111 vss 0.01873f
C704 vdd.n112 vss 0.01871f
C705 vdd.n113 vss 0.01873f
C706 vdd.n114 vss 0.11683f
C707 vdd.n115 vss 0.11683f
C708 vdd.n116 vss 0.01873f
C709 vdd.n117 vss 0.01873f
C710 vdd.n118 vss 0.01871f
C711 vdd.n119 vss 0.01873f
C712 vdd.n120 vss 0.58772f
C713 vdd.n121 vss 0.14091f
C714 vdd.n122 vss 0.58772f
C715 vdd.n123 vss 0.01873f
C716 vdd.n124 vss 0.01873f
C717 vdd.n125 vss 0.01245f
C718 vdd.n126 vss 0.01203f
C719 vdd.n127 vss 0.01263f
C720 vdd.n128 vss 0.01263f
C721 vdd.n129 vss 0.01203f
C722 vdd.n130 vss 0.00572f
C723 vdd.n131 vss 0.14091f
C724 vdd.n132 vss 0.00572f
C725 vdd.n133 vss 0.01203f
C726 vdd.n134 vss 0.01245f
C727 vdd.n135 vss 0.14091f
C728 vdd.n136 vss 0.01919f
C729 vdd.n137 vss 0.01919f
C730 vdd.n138 vss 0.00961f
C731 vdd.n139 vss 0.0067f
C732 vdd.n140 vss 0.15437f
C733 vdd.n141 vss 0.01919f
C734 vdd.n142 vss 0.01919f
C735 vdd.n143 vss 0.00961f
C736 vdd.n144 vss 0.05357f
C737 vdd.n145 vss 0.08965f
C738 vdd.n146 vss 0.08965f
C739 vdd.n147 vss 0.05327f
C740 vdd.n148 vss 0.0067f
C741 vdd.n150 vss 0.12299f
C742 vdd.n151 vss 0.01871f
C743 vdd.n152 vss 0.01873f
C744 vdd.n153 vss 0.01873f
C745 vdd.n154 vss 0.11683f
C746 vdd.n155 vss 0.11683f
C747 vdd.n156 vss 0.01873f
C748 vdd.n157 vss 0.01871f
C749 vdd.n158 vss 0.01873f
C750 vdd.n159 vss 0.01873f
C751 vdd.n160 vss 0.11772f
C752 vdd.n161 vss 0.11772f
C753 vdd.n162 vss 0.14091f
C754 vdd.n163 vss 0.01245f
C755 vdd.n164 vss 0.01245f
C756 vdd.n165 vss 0.01201f
C757 vdd.n166 vss 0.00286f
C758 vdd.n167 vss 0.14945f
C759 vdd.n168 vss 0.55066f
C760 vdd.n169 vss 0.94451f
C761 vdd.n170 vss 0.00286f
C762 vdd.n171 vss 0.16789f
C763 vdd.n172 vss 0.00288f
C764 vdd.n173 vss 0.01263f
C765 vdd.n174 vss 0.01873f
C766 vdd.n175 vss 0.01203f
C767 vdd.n176 vss 0.01873f
C768 vdd.n177 vss 0.28182f
C769 vdd.n178 vss 0.01245f
C770 vdd.n179 vss 0.01873f
C771 vdd.n180 vss 0.28182f
C772 vdd.n181 vss 0.01919f
C773 vdd.n182 vss 0.01919f
C774 vdd.n183 vss 0.01871f
C775 vdd.n184 vss 0.0067f
C776 vdd.n185 vss 0.0067f
C777 vdd.n186 vss 0.13326f
C778 vdd.n187 vss 0.00961f
C779 vdd.n188 vss 0.01919f
C780 vdd.n189 vss 0.01919f
C781 vdd.n190 vss 0.28182f
C782 vdd.n191 vss 0.01919f
C783 vdd.n192 vss 0.01919f
C784 vdd.n193 vss 0.00961f
C785 vdd.n194 vss 0.01919f
C786 vdd.n195 vss 0.01919f
C787 vdd.n196 vss 0.00961f
C788 vdd.n197 vss 0.01873f
C789 vdd.n198 vss 0.01871f
C790 vdd.n199 vss 0.01873f
C791 vdd.n200 vss 0.01873f
C792 vdd.n201 vss 0.23366f
C793 vdd.n202 vss 0.01873f
C794 vdd.n203 vss 0.01873f
C795 vdd.n204 vss 0.23366f
C796 vdd.n205 vss 0.01873f
C797 vdd.n206 vss 0.01873f
C798 vdd.n207 vss 0.01871f
C799 vdd.n208 vss 0.01873f
C800 vdd.n209 vss 0.23544f
C801 vdd.n210 vss 0.01873f
C802 vdd.n211 vss 0.01871f
C803 vdd.n212 vss 0.0067f
C804 vdd.n213 vss 0.0298f
C805 vdd.n214 vss 0.13326f
C806 vdd.n215 vss 0.02997f
C807 vdd.n216 vss 0.0067f
C808 vdd.n217 vss 0.00961f
C809 vdd.n218 vss 0.01873f
C810 vdd.n219 vss 0.01873f
C811 vdd.n220 vss 0.23544f
C812 vdd.n221 vss 0.23544f
C813 vdd.n222 vss 0.01245f
C814 vdd.n223 vss 0.01263f
C815 vdd.n224 vss 0.01203f
C816 vdd.n225 vss 0.01203f
C817 vdd.n226 vss 0.01203f
C818 vdd.n227 vss 0.28182f
C819 vdd.n228 vss 0.00572f
C820 vdd.n229 vss 0.00572f
C821 vdd.n230 vss 0.01203f
C822 vdd.n231 vss 0.01203f
C823 vdd.n232 vss 0.01245f
C824 vdd.n233 vss 0.01203f
C825 vdd.n234 vss 0.01263f
C826 vdd.n235 vss 0.01263f
C827 vdd.n236 vss 0.01201f
C828 vdd.n237 vss 0.01245f
C829 vdd.n238 vss 0.01873f
C830 vdd.n239 vss 0.01873f
C831 vdd.n240 vss 0.01203f
C832 vdd.n241 vss 0.01203f
C833 vdd.n242 vss 0.01873f
C834 vdd.n243 vss 0.01873f
C835 vdd.n244 vss 0.28182f
C836 vdd.n245 vss 0.01245f
C837 vdd.n246 vss 0.01245f
C838 vdd.n247 vss 0.01263f
C839 vdd.n248 vss 0.00288f
C840 vdd.n249 vss 0.0067f
C841 vdd.n250 vss 0.00961f
C842 vdd.n251 vss 0.01919f
C843 vdd.n252 vss 0.01919f
C844 vdd.n253 vss 0.28182f
C845 vdd.n254 vss 0.01919f
C846 vdd.n255 vss 0.01919f
C847 vdd.n256 vss 0.00961f
C848 vdd.n257 vss 0.28182f
C849 vdd.n258 vss 0.01873f
C850 vdd.n259 vss 0.01919f
C851 vdd.n260 vss 0.01919f
C852 vdd.n261 vss 0.0067f
C853 vdd.n262 vss 0.00961f
C854 vdd.n263 vss 0.01919f
C855 vdd.n264 vss 0.01919f
C856 vdd.n265 vss 0.01871f
C857 vdd.n266 vss 0.13326f
C858 vdd.n267 vss 0.04802f
C859 vdd.n268 vss 0.0067f
C860 vdd.n269 vss 0.00961f
C861 vdd.n270 vss 0.01873f
C862 vdd.n271 vss 0.01873f
C863 vdd.n272 vss 0.23544f
C864 vdd.n273 vss 0.01873f
C865 vdd.n274 vss 0.01873f
C866 vdd.n275 vss 0.01871f
C867 vdd.n276 vss 0.01873f
C868 vdd.n277 vss 0.23366f
C869 vdd.n278 vss 0.01873f
C870 vdd.n279 vss 0.01873f
C871 vdd.n280 vss 0.23366f
C872 vdd.n281 vss 0.01873f
C873 vdd.n282 vss 0.01873f
C874 vdd.n283 vss 0.01871f
C875 vdd.n284 vss 0.01873f
C876 vdd.n285 vss 0.28182f
C877 vdd.n286 vss 0.01245f
C878 vdd.n287 vss 0.01245f
C879 vdd.n288 vss 0.01203f
C880 vdd.n289 vss 0.01203f
C881 vdd.n290 vss 0.01203f
C882 vdd.n291 vss 0.00572f
C883 vdd.n292 vss 0.28182f
C884 vdd.n293 vss 0.01203f
C885 vdd.n294 vss 0.01263f
C886 vdd.n295 vss 0.01203f
C887 vdd.n296 vss 0.01203f
C888 vdd.n297 vss 0.00572f
C889 vdd.n298 vss 0.28182f
C890 vdd.n299 vss 0.28182f
C891 vdd.n300 vss 0.01263f
C892 vdd.n301 vss 0.01263f
C893 vdd.n302 vss 0.01203f
C894 vdd.n303 vss 0.01245f
C895 vdd.n304 vss 0.01873f
C896 vdd.n305 vss 0.01873f
C897 vdd.n306 vss 0.23544f
C898 vdd.n307 vss 0.23544f
C899 vdd.n308 vss 0.01873f
C900 vdd.n309 vss 0.01871f
C901 vdd.n310 vss 0.0067f
C902 vdd.n311 vss 0.0298f
C903 vdd.n312 vss 0.13326f
C904 vdd.n313 vss 0.10634f
C905 vdd.n314 vss 0.0842f
C906 vdd.n315 vss 0.00286f
C907 vdd.n316 vss 0.01201f
C908 vdd.n317 vss 0.01245f
C909 vdd.n318 vss 0.01873f
C910 vdd.n319 vss 0.01873f
C911 vdd.n320 vss 0.23544f
C912 vdd.n321 vss 0.23544f
C913 vdd.n322 vss 0.01245f
C914 vdd.n323 vss 0.01245f
C915 vdd.n324 vss 0.01873f
C916 vdd.n325 vss 0.01203f
C917 vdd.n326 vss 0.01263f
C918 vdd.n327 vss 0.01263f
C919 vdd.n328 vss 0.01203f
C920 vdd.n329 vss 0.01245f
C921 vdd.n330 vss 0.01873f
C922 vdd.n331 vss 0.01245f
C923 vdd.n332 vss 0.28182f
C924 vdd.n333 vss 0.01245f
C925 vdd.n334 vss 0.01203f
C926 vdd.n335 vss 0.01263f
C927 vdd.n336 vss 0.01263f
C928 vdd.n337 vss 0.01203f
C929 vdd.n338 vss 0.00288f
C930 vdd.n339 vss 0.00572f
C931 vdd.n340 vss 0.28182f
C932 vdd.n341 vss 0.00572f
C933 vdd.n342 vss 0.01203f
C934 vdd.n343 vss 0.01245f
C935 vdd.n344 vss 0.28182f
C936 vdd.n345 vss 0.01245f
C937 vdd.n346 vss 0.01245f
C938 vdd.n347 vss 0.01201f
C939 vdd.n348 vss 0.00286f
C940 vdd.n349 vss 0.08395f
C941 vdd.n350 vss 0.04495f
C942 vdd.n351 vss 0.61182f
C943 vdd.n352 vss 2.80783f
C944 vdd.n353 vss 0.0067f
C945 vdd.n354 vss 0.13326f
C946 vdd.n355 vss 0.00961f
C947 vdd.n356 vss 0.01919f
C948 vdd.n357 vss 0.01919f
C949 vdd.n358 vss 0.9524f
C950 vdd.n359 vss 0.01873f
C951 vdd.n360 vss 0.9524f
C952 vdd.n361 vss 0.01873f
C953 vdd.n362 vss 0.01873f
C954 vdd.n363 vss 0.01919f
C955 vdd.n364 vss 0.01919f
C956 vdd.n365 vss 0.01871f
C957 vdd.n366 vss 0.00961f
C958 vdd.n367 vss 0.01919f
C959 vdd.n368 vss 0.01919f
C960 vdd.n369 vss 0.9524f
C961 vdd.n370 vss 0.01873f
C962 vdd.n371 vss 0.01873f
C963 vdd.n372 vss 0.01873f
C964 vdd.n373 vss 0.9524f
C965 vdd.n374 vss 0.01919f
C966 vdd.n375 vss 0.01919f
C967 vdd.n376 vss 0.00961f
C968 vdd.n377 vss 0.01873f
C969 vdd.n378 vss 0.01871f
C970 vdd.n379 vss 0.01873f
C971 vdd.n380 vss 1.47703f
C972 vdd.n381 vss 0.01873f
C973 vdd.n382 vss 0.01871f
C974 vdd.n383 vss 0.0067f
C975 vdd.n384 vss 0.13326f
C976 vdd.n385 vss 0.0298f
C977 vdd.n386 vss 0.0067f
C978 vdd.n387 vss 0.00961f
C979 vdd.n388 vss 0.01873f
C980 vdd.n389 vss 0.01873f
C981 vdd.n390 vss 1.47703f
C982 vdd.n391 vss 0.01873f
C983 vdd.n392 vss 0.01871f
C984 vdd.n393 vss 0.0067f
C985 vdd.n394 vss 0.15064f
C986 vdd.n395 vss 0.81864f
C987 vdd.n396 vss 1.73787f
C988 vdd.n397 vss 0.0067f
C989 vdd.n398 vss 0.13326f
C990 vdd.n399 vss 0.00961f
C991 vdd.n400 vss 0.01919f
C992 vdd.n401 vss 0.01919f
C993 vdd.n402 vss 0.9524f
C994 vdd.n403 vss 0.01873f
C995 vdd.n404 vss 0.9524f
C996 vdd.n405 vss 0.01873f
C997 vdd.n406 vss 0.01873f
C998 vdd.n407 vss 0.01919f
C999 vdd.n408 vss 0.01919f
C1000 vdd.n409 vss 0.01871f
C1001 vdd.n410 vss 0.00961f
C1002 vdd.n411 vss 0.01919f
C1003 vdd.n412 vss 0.01919f
C1004 vdd.n413 vss 0.9524f
C1005 vdd.n414 vss 0.01873f
C1006 vdd.n415 vss 0.01873f
C1007 vdd.n416 vss 0.01873f
C1008 vdd.n417 vss 0.9524f
C1009 vdd.n418 vss 0.01919f
C1010 vdd.n419 vss 0.01919f
C1011 vdd.n420 vss 0.00961f
C1012 vdd.n421 vss 0.01873f
C1013 vdd.n422 vss 0.01871f
C1014 vdd.n423 vss 0.01873f
C1015 vdd.n424 vss 1.47703f
C1016 vdd.n425 vss 0.01873f
C1017 vdd.n426 vss 0.01871f
C1018 vdd.n427 vss 0.0067f
C1019 vdd.n428 vss 0.13326f
C1020 vdd.n429 vss 0.0298f
C1021 vdd.n430 vss 0.0067f
C1022 vdd.n431 vss 0.00961f
C1023 vdd.n432 vss 0.01873f
C1024 vdd.n433 vss 0.01873f
C1025 vdd.n434 vss 1.47703f
C1026 vdd.n435 vss 0.01873f
C1027 vdd.n436 vss 0.01871f
C1028 vdd.n437 vss 0.0067f
C1029 vdd.n438 vss 0.15064f
C1030 vdd.n439 vss 0.82009f
C1031 vdd.n440 vss 3.28978f
C1032 vdd.n441 vss 5.20077f
C1033 vdd.n442 vss 2.5442f
C1034 vdd.n443 vss 0.54218f
C1035 vdd.n444 vss 0.01748f
C1036 vdd.n445 vss 0.44609f
C1037 vdd.n446 vss 0.48123f
C1038 vdd.n447 vss 0.02158f
C1039 vdd.n448 vss 0.25936f
C1040 vdd.n449 vss 0.03904f
C1041 vdd.n450 vss 0.04413f
C1042 vdd.n451 vss 2.75905f
C1043 vdd.n452 vss 0.03916f
C1044 vdd.n453 vss 0.03916f
C1045 vdd.n454 vss 0.49708f
C1046 vdd.n455 vss 0.03904f
C1047 vdd.n456 vss 0.04413f
C1048 vdd.n457 vss 0.14251f
C1049 vdd.n458 vss -0.10005f
C1050 vdd.n459 vss 0.02158f
C1051 vdd.n460 vss 0.04413f
C1052 vdd.n461 vss 0.03615f
C1053 vdd.n462 vss 0.61995f
C1054 vdd.n463 vss 0.03916f
C1055 vdd.n464 vss 2.69761f
C1056 vdd.n465 vss 0.03916f
C1057 vdd.n466 vss 0.13183f
C1058 vdd.n467 vss 0.25716f
C1059 vdd.n468 vss 0.81131f
C1060 vdd.n469 vss 0.05057f
C1061 vdd.n470 vss 0.05057f
C1062 vdd.n471 vss 3.02434f
C1063 vdd.n472 vss 0.05057f
C1064 vdd.n473 vss 0.05057f
C1065 vdd.n474 vss 0.03615f
C1066 vdd.n475 vss 0.04413f
C1067 vdd.n476 vss 0.25716f
C1068 vdd.n477 vss 0.81131f
C1069 vdd.n478 vss 0.13183f
C1070 vdd.n479 vss 0.13091f
C1071 vdd.n480 vss 0.14124f
C1072 vdd.n481 vss 0.45695f
C1073 vdd.n482 vss 0.05028f
C1074 vdd.n483 vss 0.05047f
C1075 vdd.n484 vss 0.83064f
C1076 vdd.n485 vss 0.27172f
C1077 vdd.n486 vss 3.15001f
C1078 vdd.n487 vss 0.06016f
C1079 vdd.n488 vss 3.02434f
C1080 vdd.n489 vss 0.05045f
C1081 vdd.n490 vss 0.05045f
C1082 vdd.n491 vss 0.81131f
C1083 vdd.n492 vss 0.01835f
C1084 vdd.n493 vss 0.27172f
C1085 vdd.n494 vss 0.05028f
C1086 vdd.n495 vss 0.06041f
C1087 vdd.n496 vss 3.16397f
C1088 vdd.n497 vss 0.05047f
C1089 vdd.n498 vss 0.05047f
C1090 vdd.n499 vss 2.23126f
C1091 vdd.n500 vss 0.05028f
C1092 vdd.n501 vss 0.06041f
C1093 vdd.n502 vss 0.05028f
C1094 vdd.n503 vss 0.25936f
C1095 vdd.n504 vss 0.00715f
C1096 vdd.n505 vss 0.05057f
C1097 vdd.n506 vss 0.0514f
C1098 vdd.n507 vss -0.10005f
C1099 vdd.n508 vss 3.11929f
C1100 vdd.n509 vss 0.05057f
C1101 vdd.n510 vss 0.05028f
C1102 vdd.n511 vss 0.01835f
C1103 vdd.n512 vss 2.75905f
C1104 vdd.n513 vss 0.0514f
C1105 vdd.n514 vss 0.0514f
C1106 vdd.n515 vss 0.13743f
C1107 vdd.n516 vss 0.13118f
C1108 vdd.n517 vss 0.02158f
C1109 vdd.n518 vss 0.03904f
C1110 vdd.n519 vss 0.03916f
C1111 vdd.n520 vss 0.03615f
C1112 vdd.n521 vss 0.25716f
C1113 vdd.n522 vss 0.04413f
C1114 vdd.n523 vss 0.03916f
C1115 vdd.n524 vss 0.03916f
C1116 vdd.n525 vss 0.44293f
C1117 vdd.n526 vss 0.02369f
C1118 vdd.n527 vss 0.13183f
C1119 vdd.n528 vss 0.13091f
C1120 vdd.n529 vss 0.14124f
C1121 vdd.n530 vss 0.14251f
C1122 vdd.n531 vss 0.00715f
C1123 vdd.n532 vss 0.45695f
C1124 vdd.n533 vss 0.83064f
C1125 vdd.n534 vss 0.25936f
C1126 vdd.n535 vss 2.56357f
C1127 vdd.n536 vss 0.03916f
C1128 vdd.n537 vss 0.03904f
C1129 vdd.n538 vss 0.03615f
C1130 vdd.n539 vss 0.12816f
C1131 vdd.n540 vss 0.03916f
C1132 vdd.n541 vss 0.04413f
C1133 vdd.n542 vss 0.13183f
C1134 vdd.n543 vss 2.2145f
C1135 vdd.n544 vss 0.13091f
C1136 vdd.n545 vss 0.13118f
C1137 vdd.n546 vss 0.14251f
C1138 vdd.n547 vss 0.14124f
C1139 vdd.n548 vss 0.01835f
C1140 vdd.n549 vss 0.01835f
C1141 vdd.n550 vss 0.05028f
C1142 vdd.n551 vss 0.05045f
C1143 vdd.n552 vss 0.61995f
C1144 vdd.n553 vss 0.05045f
C1145 vdd.n554 vss 0.04638f
C1146 vdd.n555 vss 0.27022f
C1147 vdd.n556 vss 0.25716f
C1148 vdd.n557 vss 0.81131f
C1149 vdd.n558 vss 0.44293f
C1150 vdd.n559 vss 0.02369f
C1151 vdd.n560 vss 0.13743f
C1152 vdd.n561 vss 0.03916f
C1153 vdd.n562 vss 0.03904f
C1154 vdd.n563 vss 0.00818f
C1155 vdd.n564 vss 0.00818f
C1156 vdd.n565 vss 0.02158f
C1157 vdd.n566 vss 0.83837f
C1158 vdd.n567 vss 0.0361f
C1159 vdd.n568 vss 0.01748f
C1160 vdd.n569 vss 0.63588f
C1161 vdd.n570 vss 0.21788f
C1162 vdd.n571 vss 1.9946f
C1163 vdd.n572 vss 0.72756f
C1164 vdd.n573 vss 0.72296f
C1165 vdd.n574 vss 0.02158f
C1166 vdd.n575 vss 0.25936f
C1167 vdd.n576 vss 0.03904f
C1168 vdd.n577 vss 0.04413f
C1169 vdd.n578 vss 1.37952f
C1170 vdd.n579 vss 0.03916f
C1171 vdd.n580 vss 0.05047f
C1172 vdd.n581 vss 1.11563f
C1173 vdd.n582 vss 0.05028f
C1174 vdd.n583 vss 1.575f
C1175 vdd.n584 vss 0.90878f
C1176 vdd.n585 vss 0.05057f
C1177 vdd.n586 vss 0.05057f
C1178 vdd.n587 vss 0.05058f
C1179 vdd.n589 vss 0.5841f
C1180 vdd.n590 vss 0.02893f
C1181 vdd.n591 vss 0.80452f
C1182 vdd.n592 vss 0.36147f
C1183 vdd.n593 vss 0.23958f
C1184 vdd.n594 vss 0.23624f
C1185 vdd.n595 vss 0.02863f
C1186 vdd.n596 vss 0.05279f
C1187 vdd.n597 vss 0.0514f
C1188 vdd.n598 vss 1.43378f
C1189 vdd.n599 vss 2.1583f
C1190 vdd.n600 vss 0.06041f
C1191 vdd.n601 vss 0.14251f
C1192 vdd.n602 vss 0.83064f
C1193 vdd.n603 vss 0.05057f
C1194 vdd.n604 vss 0.0514f
C1195 vdd.n605 vss -0.10005f
C1196 vdd.n606 vss 0.30997f
C1197 vdd.n607 vss 0.13118f
C1198 vdd.n608 vss 0.12816f
C1199 vdd.n609 vss 0.00818f
C1200 vdd.n610 vss 0.00818f
C1201 vdd.n611 vss 0.03904f
C1202 vdd.n612 vss 0.03916f
C1203 vdd.n613 vss 0.04413f
C1204 vdd.n614 vss 0.27022f
C1205 vdd.n615 vss 0.13091f
C1206 vdd.n616 vss 0.05028f
C1207 vdd.n617 vss 0.14124f
C1208 vdd.n618 vss 0.01835f
C1209 vdd.n619 vss 0.01835f
C1210 vdd.n620 vss 0.27172f
C1211 vdd.n621 vss 0.04637f
C1212 vdd.n622 vss 0.05028f
C1213 vdd.n623 vss 0.04638f
C1214 vdd.n624 vss 0.05045f
C1215 vdd.n625 vss 1.10725f
C1216 vdd.n626 vss 1.6455f
C1217 vdd.n627 vss 1.21001f
C1218 vdd.n628 vss 0.05045f
C1219 vdd.n629 vss 0.13183f
C1220 vdd.n630 vss 0.13743f
C1221 vdd.n631 vss 0.02369f
C1222 vdd.n632 vss 0.44293f
C1223 vdd.n633 vss 0.81131f
C1224 vdd.n634 vss 0.25716f
C1225 vdd.n635 vss 0.03615f
C1226 vdd.n636 vss 0.03916f
C1227 vdd.n637 vss 1.55964f
C1228 vdd.n638 vss 1.34881f
C1229 vdd.n639 vss 0.05057f
C1230 vdd.n640 vss 0.0514f
C1231 vdd.n641 vss 0.45695f
C1232 vdd.n642 vss 0.00715f
C1233 vdd.n643 vss 0.05047f
C1234 vdd.n644 vss 0.24854f
C1235 vdd.n645 vss 1.58198f
C1236 vdd.n646 vss 0.03916f
C1237 vdd.n647 vss 0.0361f
C1238 vdd.n648 vss 0.01748f
C1239 vdd.n649 vss 0.03864f
C1240 vdd.n650 vss 0.52001f
C1241 vdd.n651 vss 0.39387f
C1242 vdd.n652 vss 0.33632f
C1243 vdd.n653 vss 1.25631f
C1244 vdd.n654 vss 4.49433f
C1245 vdd.n655 vss 2.68756f
C1246 vdd.n656 vss 0.22801f
C1247 vdd.n657 vss 3.71924f
C1248 vdd.n658 vss 0.09907f
C1249 vdd.n659 vss 0.44609f
C1250 vdd.n660 vss 0.48123f
C1251 vdd.n661 vss 0.02879f
C1252 vdd.n662 vss 0.01748f
C1253 vdd.n663 vss 0.0361f
C1254 vdd.n664 vss 0.03916f
C1255 vdd.n665 vss 0.04413f
C1256 vdd.n666 vss 3.15001f
C1257 vdd.n667 vss 0.04413f
C1258 vdd.n668 vss 0.03916f
C1259 vdd.n669 vss 0.03904f
C1260 vdd.n670 vss 0.00818f
C1261 vdd.n671 vss 0.00818f
C1262 vdd.n672 vss 0.12816f
C1263 vdd.n673 vss -0.10005f
C1264 vdd.n674 vss 0.05057f
C1265 vdd.n675 vss 2.69761f
C1266 vdd.n676 vss 0.05057f
C1267 vdd.n677 vss 0.0514f
C1268 vdd.n678 vss 0.45695f
C1269 vdd.n679 vss 0.83064f
C1270 vdd.n680 vss 0.27172f
C1271 vdd.n681 vss 0.04637f
C1272 vdd.n682 vss 0.05047f
C1273 vdd.n683 vss 0.49708f
C1274 vdd.n684 vss 0.05047f
C1275 vdd.n685 vss 0.04637f
C1276 vdd.n686 vss 0.05028f
C1277 vdd.n687 vss 0.04638f
C1278 vdd.n688 vss 0.27022f
C1279 vdd.n689 vss 0.06016f
C1280 vdd.n690 vss 3.29522f
C1281 vdd.n691 vss 0.05047f
C1282 vdd.n692 vss 0.05047f
C1283 vdd.n693 vss 0.13091f
C1284 vdd.n694 vss 0.14124f
C1285 vdd.n695 vss 0.01835f
C1286 vdd.n696 vss 0.27022f
C1287 vdd.n697 vss 0.05045f
C1288 vdd.n698 vss 0.05045f
C1289 vdd.n699 vss 0.04637f
C1290 vdd.n700 vss 0.05028f
C1291 vdd.n701 vss 0.01835f
C1292 vdd.n702 vss 0.01835f
C1293 vdd.n703 vss 0.05028f
C1294 vdd.n704 vss 0.04638f
C1295 vdd.n705 vss 0.27022f
C1296 vdd.n706 vss 0.06016f
C1297 vdd.n707 vss 2.56636f
C1298 vdd.n708 vss 0.06016f
C1299 vdd.n709 vss 0.05045f
C1300 vdd.n710 vss 0.05028f
C1301 vdd.n711 vss 0.01835f
C1302 vdd.n712 vss 0.05028f
C1303 vdd.n713 vss 0.05045f
C1304 vdd.n714 vss 0.04638f
C1305 vdd.n715 vss 0.05028f
C1306 vdd.n716 vss 0.04637f
C1307 vdd.n717 vss 0.0361f
C1308 vdd.n718 vss 0.25936f
C1309 vdd.n719 vss 0.00715f
C1310 vdd.n720 vss 0.0514f
C1311 vdd.n721 vss 2.23126f
C1312 vdd.n722 vss 0.0514f
C1313 vdd.n723 vss 0.45695f
C1314 vdd.n724 vss 0.83064f
C1315 vdd.n725 vss 0.27172f
C1316 vdd.n726 vss 0.06041f
C1317 vdd.n727 vss 3.29801f
C1318 vdd.n728 vss 0.06041f
C1319 vdd.n729 vss 0.05047f
C1320 vdd.n730 vss 0.00715f
C1321 vdd.n731 vss 0.14251f
C1322 vdd.n732 vss 0.13118f
C1323 vdd.n733 vss 0.03904f
C1324 vdd.n734 vss 0.00818f
C1325 vdd.n735 vss 0.00818f
C1326 vdd.n736 vss 0.12816f
C1327 vdd.n737 vss -0.10005f
C1328 vdd.n738 vss 0.13743f
C1329 vdd.n739 vss 0.02369f
C1330 vdd.n740 vss 0.44293f
C1331 vdd.n741 vss 0.0514f
C1332 vdd.n742 vss 2.2145f
C1333 vdd.n743 vss 0.0514f
C1334 vdd.n744 vss 0.44293f
C1335 vdd.n745 vss 0.02369f
C1336 vdd.n746 vss 0.13743f
C1337 vdd.n747 vss 0.03916f
C1338 vdd.n748 vss 3.11929f
C1339 vdd.n749 vss 0.03916f
C1340 vdd.n750 vss 0.03904f
C1341 vdd.n751 vss 0.00818f
C1342 vdd.n752 vss 0.00818f
C1343 vdd.n753 vss 0.12816f
C1344 vdd.n754 vss 0.13118f
C1345 vdd.n755 vss 0.03916f
C1346 vdd.n756 vss 3.16397f
C1347 vdd.n757 vss 0.03916f
C1348 vdd.n758 vss 0.0361f
C1349 vdd.n759 vss 0.01748f
C1350 vdd.n760 vss 0.02879f
C1351 vdd.n761 vss 0.83837f
C1352 vdd.n762 vss 0.63604f
C1353 vdd.n763 vss 4.00496f
C1354 vdd.n764 vss 13.4458f
C1355 vdd.n765 vss 2.61538f
C1356 vdd.n766 vss 2.17134f
C1357 vdd.n767 vss 0.97747f
C1358 vdd.n768 vss 0.90807f
C1359 vdd.n769 vss 0.49766f
C1360 vdd.n770 vss 0.69026f
C1361 vdd.n771 vss 0.05342f
C1362 vdd.n772 vss 0.01748f
C1363 vdd.n773 vss 0.0361f
C1364 vdd.n774 vss 0.25936f
C1365 vdd.n775 vss 0.04413f
C1366 vdd.n776 vss 0.03916f
C1367 vdd.n777 vss 0.13118f
C1368 vdd.n778 vss 0.12816f
C1369 vdd.n779 vss 0.00818f
C1370 vdd.n780 vss 0.00818f
C1371 vdd.n781 vss 1.37952f
C1372 vdd.n782 vss 0.01835f
C1373 vdd.n783 vss 0.01835f
C1374 vdd.n784 vss 0.05028f
C1375 vdd.n785 vss 0.04637f
C1376 vdd.n786 vss 0.27172f
C1377 vdd.n787 vss 0.06041f
C1378 vdd.n788 vss 1.64901f
C1379 vdd.n789 vss 1.64761f
C1380 vdd.n790 vss 1.51217f
C1381 vdd.n791 vss 0.04413f
C1382 vdd.n792 vss 0.0514f
C1383 vdd.n793 vss 0.0348f
C1384 vdd.n794 vss 0.05024f
C1385 vdd.n795 vss 1.34881f
C1386 vdd.n796 vss 0.06708f
C1387 vdd.n797 vss 0.05949f
C1388 vdd.n798 vss 0.1282f
C1389 vdd.n799 vss 0.13064f
C1390 vdd.n800 vss 0.00818f
C1391 vdd.n801 vss 0.00818f
C1392 vdd.n802 vss 0.03904f
C1393 vdd.n803 vss 0.03916f
C1394 vdd.n804 vss 0.13392f
C1395 vdd.n805 vss 0.02369f
C1396 vdd.n806 vss 0.13183f
C1397 vdd.n807 vss 0.05045f
C1398 vdd.n808 vss 0.30997f
C1399 vdd.n809 vss 0.05045f
C1400 vdd.n810 vss 0.05028f
C1401 vdd.n811 vss 0.01835f
C1402 vdd.n812 vss 0.01835f
C1403 vdd.n813 vss 0.14124f
C1404 vdd.n814 vss 0.13471f
C1405 vdd.n815 vss 0.0524f
C1406 vdd.n816 vss 0.24854f
C1407 vdd.n817 vss 1.58198f
C1408 vdd.n818 vss 0.03667f
C1409 vdd.n819 vss 0.03574f
C1410 vdd.n820 vss 0.01748f
C1411 vdd.n821 vss 0.05342f
C1412 vdd.n822 vss 0.90807f
C1413 vdd.n823 vss 0.97747f
C1414 vdd.n824 vss 2.46713f
C1415 vdd.n825 vss 0.19222f
C1416 vdd.n826 vss 0.14978f
C1417 vdd.n827 vss 0.17304f
C1418 comp_p_6/vbias_p.t3 vss 0.68603f
C1419 comp_p_6/vbias_p.t2 vss 0.72096f
C1420 comp_p_6/vbias_p.n0 vss 1.08732f
C1421 comp_p_6/vbias_p.n1 vss 1.83502f
C1422 comp_p_6/vbias_p.t4 vss 0.68603f
C1423 comp_p_6/vbias_p.t6 vss 0.68603f
C1424 comp_p_6/vbias_p.t5 vss 0.68603f
C1425 comp_p_6/vbias_p.t7 vss 0.68603f
C1426 comp_p_6/vbias_p.n2 vss 2.59376f
C1427 comp_p_6/vbias_p.n3 vss 3.00057f
C1428 comp_p_6/vbias_p.n4 vss 0.88625f
C1429 comp_p_6/vbias_p.n5 vss 9.0963f
C1430 comp_p_6/vbias_p.n6 vss 0.28438f
C1431 comp_p_6/vbias_p.t0 vss 0.66673f
C1432 comp_p_6/vbias_p.t8 vss 0.72096f
C1433 comp_p_6/vbias_p.n7 vss 0.24366f
C1434 comp_p_6/vbias_p.n8 vss 1.20496f
C1435 comp_p_6/vbias_p.t1 vss 0.26393f
C1436 tmux_7therm_to_3bin_0/tmux_2to1_3/A vss 0.4939f
C1437 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G vss 0.55051f
C1438 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin vss 0.52606f
C1439 dout2 vss 0.32356f
C1440 tmux_7therm_to_3bin_0/buffer_8/inv_1/vin vss 0.52606f
C1441 dout1 vss 0.32356f
C1442 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vss 0.52606f
C1443 dout0 vss 0.32356f
C1444 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin vss 0.52765f
C1445 tmux_7therm_to_3bin_0/buffer_6/out vss 0.67609f
C1446 d6 vss -14.33288f
C1447 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin vss 0.52606f
C1448 tmux_7therm_to_3bin_0/buffer_5/out vss 0.70857f
C1449 d5 vss 10.50535f
C1450 vdd vss 0.37121p
C1451 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vss 0.52606f
C1452 tmux_7therm_to_3bin_0/buffer_4/out vss 0.70167f
C1453 d4 vss 10.04751f
C1454 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin vss 0.52606f
C1455 tmux_7therm_to_3bin_0/R1/R2 vss 0.22083f
C1456 d3 vss 3.16422f
C1457 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin vss 0.52811f
C1458 tmux_7therm_to_3bin_0/buffer_2/out vss 0.28552f
C1459 d2 vss 7.17248f
C1460 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin vss 0.52606f
C1461 tmux_7therm_to_3bin_0/buffer_1/out vss 0.30295f
C1462 d1 vss 10.33787f
C1463 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin vss 0.52606f
C1464 tmux_7therm_to_3bin_0/buffer_0/out vss 0.30577f
C1465 d0 vss 6.01917f
C1466 tmux_7therm_to_3bin_0/R1/m1_n100_n100# vss 0.10692f
C1467 tmux_7therm_to_3bin_0/buffer_8/in vss 1.28735f
C1468 tmux_7therm_to_3bin_0/buffer_7/in vss 0.74661f
C1469 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vss 0.55051f
C1470 tmux_7therm_to_3bin_0/R1/R1 vss 3.00001f
C1471 tmux_7therm_to_3bin_0/tmux_2to1_3/B vss 0.41874f
C1472 tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G vss 0.55051f
C1473 tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G vss 0.55051f
C1474 vin vss 23.06873f
C1475 comp_p_6/tail vss 1.09633f
C1476 comp_p_6/latch_right vss 3.49411f
C1477 comp_p_6/out_left vss 3.20258f
C1478 comp_p_6/latch_left vss 10.479f
C1479 comp_p_5/tail vss 1.09613f
C1480 comp_p_5/latch_right vss 3.49805f
C1481 comp_p_5/out_left vss 2.08667f
C1482 comp_p_5/latch_left vss 10.47837f
C1483 comp_p_4/tail vss 1.56897f
C1484 comp_p_4/latch_right vss 5.50989f
C1485 comp_p_4/out_left vss 5.17613f
C1486 comp_p_4/latch_left vss 11.51511f
C1487 comp_p_3/tail vss 1.09611f
C1488 comp_p_3/latch_right vss 12.24146f
C1489 comp_p_3/out_left vss 3.17448f
C1490 comp_p_3/latch_left vss 10.47733f
C1491 comp_p_2/tail vss 1.56898f
C1492 comp_p_2/latch_right vss 5.49653f
C1493 comp_p_2/out_left vss 4.34035f
C1494 comp_p_2/latch_left vss 11.51222f
C1495 comp_p_0/tail vss 1.56897f
C1496 comp_p_0/latch_right vss 5.50255f
C1497 comp_p_0/out_left vss 5.23512f
C1498 comp_p_0/latch_left vss 6.03535f
C1499 comp_p_1/tail vss 1.09611f
C1500 comp_p_1/latch_right vss 3.49227f
C1501 comp_p_1/out_left vss 2.0627f
C1502 comp_p_1/latch_left vss 10.47733f
C1503 comp_p_0/vinn vss 6.06348f
C1504 comp_p_2/vinn vss 4.46291f
C1505 comp_p_3/vinn vss 7.47636f
C1506 comp_p_4/vinn vss 4.49649f
C1507 comp_p_5/vinn vss 7.17599f
C1508 comp_p_6/vinn vss 8.16656f
C1509 comp_p_1/vinn vss 8.18212f
C1510 vref vss 4.52985f
C1511 vbias_generation_0/bias_n vss 2.63421f
C1512 vbias_generation_0/XR_bias_4/R1 vss 1.61917f
C1513 vbias_generation_0/XR_bias_3/R2 vss 1.9113f
C1514 vbias_generation_0/XR_bias_2/R2 vss 1.5274f
C1515 comp_p_6/vbias_p vss 22.45594f
.ends

