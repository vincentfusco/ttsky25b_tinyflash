VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tinyflash
  CLASS BLOCK ;
  FOREIGN tt_um_tinyflash ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 60.560 146.290 72.110 215.420 ;
      LAYER nwell ;
        RECT 73.730 202.210 126.150 215.330 ;
      LAYER pwell ;
        RECT 73.730 191.430 126.150 202.210 ;
      LAYER nwell ;
        RECT 73.730 165.190 126.150 191.430 ;
      LAYER pwell ;
        RECT 73.730 159.800 126.150 165.190 ;
      LAYER nwell ;
        RECT 127.890 210.860 146.850 215.050 ;
      LAYER pwell ;
        RECT 127.890 204.660 146.850 210.860 ;
      LAYER nwell ;
        RECT 127.890 196.280 146.850 204.660 ;
      LAYER pwell ;
        RECT 127.890 193.180 146.850 196.280 ;
        RECT 127.890 192.890 143.380 193.180 ;
        RECT 145.630 192.890 146.850 193.180 ;
        RECT 127.890 190.080 146.850 192.890 ;
      LAYER nwell ;
        RECT 127.890 181.700 146.850 190.080 ;
      LAYER pwell ;
        RECT 127.890 175.500 146.850 181.700 ;
      LAYER nwell ;
        RECT 127.890 167.120 146.850 175.500 ;
      LAYER pwell ;
        RECT 127.890 164.020 146.850 167.120 ;
        RECT 100.530 154.410 126.140 159.800 ;
        RECT 84.010 141.590 97.570 154.410 ;
      LAYER nwell ;
        RECT 97.570 141.590 126.140 154.410 ;
        RECT 100.530 141.290 126.140 141.590 ;
      LAYER li1 ;
        RECT 60.740 215.070 71.930 215.240 ;
        RECT 60.740 208.380 60.910 215.070 ;
        RECT 61.390 208.860 63.550 214.590 ;
        RECT 69.120 208.860 71.280 214.590 ;
        RECT 71.760 208.380 71.930 215.070 ;
        RECT 60.740 208.210 71.930 208.380 ;
        RECT 60.740 201.520 60.910 208.210 ;
        RECT 61.390 202.000 63.550 207.730 ;
        RECT 69.120 202.000 71.280 207.730 ;
        RECT 71.760 201.520 71.930 208.210 ;
        RECT 73.900 214.980 99.160 215.150 ;
        RECT 73.900 212.720 76.970 214.980 ;
        RECT 77.685 214.410 85.725 214.580 ;
        RECT 77.300 213.350 77.470 214.350 ;
        RECT 85.940 213.350 86.110 214.350 ;
        RECT 77.685 213.120 85.725 213.290 ;
        RECT 86.450 212.720 86.620 214.980 ;
        RECT 87.345 214.410 95.385 214.580 ;
        RECT 86.960 213.350 87.130 214.350 ;
        RECT 95.600 213.350 95.770 214.350 ;
        RECT 87.345 213.120 95.385 213.290 ;
        RECT 96.110 212.730 99.160 214.980 ;
        RECT 92.380 212.720 99.160 212.730 ;
        RECT 73.900 212.110 99.160 212.720 ;
        RECT 73.900 209.850 80.900 212.110 ;
        RECT 81.705 211.710 91.585 212.110 ;
        RECT 81.625 211.540 91.665 211.710 ;
        RECT 81.240 210.480 81.410 211.480 ;
        RECT 91.880 210.480 92.050 211.480 ;
        RECT 81.625 210.250 91.665 210.420 ;
        RECT 92.380 209.850 99.160 212.110 ;
        RECT 73.900 208.770 99.160 209.850 ;
        RECT 73.900 203.700 75.260 208.770 ;
        RECT 75.835 208.270 85.870 208.440 ;
        RECT 75.450 207.860 75.620 208.210 ;
        RECT 86.085 207.860 86.255 208.210 ;
        RECT 75.835 207.630 85.870 207.800 ;
        RECT 75.835 207.070 85.870 207.240 ;
        RECT 75.450 206.660 75.620 207.010 ;
        RECT 86.085 206.660 86.255 207.010 ;
        RECT 75.835 206.430 85.870 206.600 ;
        RECT 75.835 205.870 85.870 206.040 ;
        RECT 75.450 205.460 75.620 205.810 ;
        RECT 86.085 205.460 86.255 205.810 ;
        RECT 75.835 205.230 85.870 205.400 ;
        RECT 75.835 204.670 85.870 204.840 ;
        RECT 75.450 204.260 75.620 204.610 ;
        RECT 86.085 204.260 86.255 204.610 ;
        RECT 75.835 204.030 85.870 204.200 ;
        RECT 86.450 203.700 86.620 208.770 ;
        RECT 87.195 208.270 97.230 208.440 ;
        RECT 86.810 207.860 86.980 208.210 ;
        RECT 96.470 207.800 97.190 207.880 ;
        RECT 97.445 207.860 97.615 208.210 ;
        RECT 87.195 207.630 97.230 207.800 ;
        RECT 96.470 207.540 97.190 207.630 ;
        RECT 87.195 207.070 97.230 207.240 ;
        RECT 86.810 206.660 86.980 207.010 ;
        RECT 97.445 206.660 97.615 207.010 ;
        RECT 87.195 206.430 97.230 206.600 ;
        RECT 87.195 205.870 97.230 206.040 ;
        RECT 86.810 205.460 86.980 205.810 ;
        RECT 96.470 205.400 97.190 205.480 ;
        RECT 97.445 205.460 97.615 205.810 ;
        RECT 87.195 205.230 97.230 205.400 ;
        RECT 96.470 205.140 97.190 205.230 ;
        RECT 87.195 204.670 97.230 204.840 ;
        RECT 86.810 204.260 86.980 204.610 ;
        RECT 97.445 204.260 97.615 204.610 ;
        RECT 87.195 204.030 97.230 204.200 ;
        RECT 97.805 203.700 99.160 208.770 ;
        RECT 73.900 203.530 99.160 203.700 ;
        RECT 100.710 214.980 125.970 215.150 ;
        RECT 100.710 212.720 103.780 214.980 ;
        RECT 104.495 214.410 112.535 214.580 ;
        RECT 104.110 213.350 104.280 214.350 ;
        RECT 112.750 213.350 112.920 214.350 ;
        RECT 104.495 213.120 112.535 213.290 ;
        RECT 113.260 212.720 113.430 214.980 ;
        RECT 114.155 214.410 122.195 214.580 ;
        RECT 113.770 213.350 113.940 214.350 ;
        RECT 122.410 213.350 122.580 214.350 ;
        RECT 114.155 213.120 122.195 213.290 ;
        RECT 122.920 212.730 125.970 214.980 ;
        RECT 128.090 214.870 129.790 214.910 ;
        RECT 130.190 214.870 131.890 214.910 ;
        RECT 142.840 214.870 144.540 214.910 ;
        RECT 144.940 214.870 146.640 214.910 ;
        RECT 119.190 212.720 125.970 212.730 ;
        RECT 100.710 212.110 125.970 212.720 ;
        RECT 100.710 209.850 107.710 212.110 ;
        RECT 108.515 211.710 118.395 212.110 ;
        RECT 108.435 211.540 118.475 211.710 ;
        RECT 108.050 210.480 108.220 211.480 ;
        RECT 118.690 210.480 118.860 211.480 ;
        RECT 108.435 210.250 118.475 210.420 ;
        RECT 119.190 209.850 125.970 212.110 ;
        RECT 128.070 214.700 129.820 214.870 ;
        RECT 128.070 211.210 128.240 214.700 ;
        RECT 128.780 214.190 129.110 214.360 ;
        RECT 128.640 211.935 128.810 213.975 ;
        RECT 129.080 211.935 129.250 213.975 ;
        RECT 128.780 211.550 129.110 211.720 ;
        RECT 129.650 211.210 129.820 214.700 ;
        RECT 128.070 211.040 129.820 211.210 ;
        RECT 130.170 214.700 131.920 214.870 ;
        RECT 130.170 211.210 130.340 214.700 ;
        RECT 130.880 214.190 131.210 214.360 ;
        RECT 130.740 211.935 130.910 213.975 ;
        RECT 131.180 211.935 131.350 213.975 ;
        RECT 130.880 211.550 131.210 211.720 ;
        RECT 131.750 211.210 131.920 214.700 ;
        RECT 130.170 211.040 131.920 211.210 ;
        RECT 132.280 214.700 137.190 214.870 ;
        RECT 132.280 211.210 132.450 214.700 ;
        RECT 132.990 214.190 133.320 214.360 ;
        RECT 132.850 211.935 133.020 213.975 ;
        RECT 133.290 211.935 133.460 213.975 ;
        RECT 132.990 211.550 133.320 211.720 ;
        RECT 133.860 211.210 134.030 214.700 ;
        RECT 134.570 214.190 134.900 214.360 ;
        RECT 134.430 211.935 134.600 213.975 ;
        RECT 134.870 211.935 135.040 213.975 ;
        RECT 134.570 211.550 134.900 211.720 ;
        RECT 135.440 211.210 135.610 214.700 ;
        RECT 136.150 214.190 136.480 214.360 ;
        RECT 136.010 211.935 136.180 213.975 ;
        RECT 136.450 211.935 136.620 213.975 ;
        RECT 136.150 211.550 136.480 211.720 ;
        RECT 137.020 211.210 137.190 214.700 ;
        RECT 132.280 211.040 137.190 211.210 ;
        RECT 142.820 214.700 144.570 214.870 ;
        RECT 142.820 211.210 142.990 214.700 ;
        RECT 143.530 214.190 143.860 214.360 ;
        RECT 143.390 211.935 143.560 213.975 ;
        RECT 143.830 211.935 144.000 213.975 ;
        RECT 143.530 211.550 143.860 211.720 ;
        RECT 144.400 211.210 144.570 214.700 ;
        RECT 142.820 211.040 144.570 211.210 ;
        RECT 144.920 214.700 146.670 214.870 ;
        RECT 144.920 211.210 145.090 214.700 ;
        RECT 145.630 214.190 145.960 214.360 ;
        RECT 145.490 211.935 145.660 213.975 ;
        RECT 145.930 211.935 146.100 213.975 ;
        RECT 145.630 211.550 145.960 211.720 ;
        RECT 146.500 211.210 146.670 214.700 ;
        RECT 144.920 211.040 146.670 211.210 ;
        RECT 100.710 208.770 125.970 209.850 ;
        RECT 100.710 203.700 102.070 208.770 ;
        RECT 102.645 208.270 112.680 208.440 ;
        RECT 102.260 207.860 102.430 208.210 ;
        RECT 112.895 207.860 113.065 208.210 ;
        RECT 102.645 207.630 112.680 207.800 ;
        RECT 102.645 207.070 112.680 207.240 ;
        RECT 102.260 206.660 102.430 207.010 ;
        RECT 112.895 206.660 113.065 207.010 ;
        RECT 102.645 206.430 112.680 206.600 ;
        RECT 102.645 205.870 112.680 206.040 ;
        RECT 102.260 205.460 102.430 205.810 ;
        RECT 112.895 205.460 113.065 205.810 ;
        RECT 102.645 205.230 112.680 205.400 ;
        RECT 102.645 204.670 112.680 204.840 ;
        RECT 102.260 204.260 102.430 204.610 ;
        RECT 112.895 204.260 113.065 204.610 ;
        RECT 102.645 204.030 112.680 204.200 ;
        RECT 113.260 203.700 113.430 208.770 ;
        RECT 114.005 208.270 124.040 208.440 ;
        RECT 113.620 207.860 113.790 208.210 ;
        RECT 123.280 207.800 124.000 207.880 ;
        RECT 124.255 207.860 124.425 208.210 ;
        RECT 114.005 207.630 124.040 207.800 ;
        RECT 123.280 207.540 124.000 207.630 ;
        RECT 114.005 207.070 124.040 207.240 ;
        RECT 113.620 206.660 113.790 207.010 ;
        RECT 124.255 206.660 124.425 207.010 ;
        RECT 114.005 206.430 124.040 206.600 ;
        RECT 114.005 205.870 124.040 206.040 ;
        RECT 113.620 205.460 113.790 205.810 ;
        RECT 123.280 205.400 124.000 205.480 ;
        RECT 124.255 205.460 124.425 205.810 ;
        RECT 114.005 205.230 124.040 205.400 ;
        RECT 123.280 205.140 124.000 205.230 ;
        RECT 114.005 204.670 124.040 204.840 ;
        RECT 113.620 204.260 113.790 204.610 ;
        RECT 124.255 204.260 124.425 204.610 ;
        RECT 114.005 204.030 124.040 204.200 ;
        RECT 124.615 203.700 125.970 208.770 ;
        RECT 128.070 210.510 129.820 210.680 ;
        RECT 128.070 208.110 128.240 210.510 ;
        RECT 128.780 210.000 129.110 210.170 ;
        RECT 128.640 208.790 128.810 209.830 ;
        RECT 129.080 208.790 129.250 209.830 ;
        RECT 128.780 208.450 129.110 208.620 ;
        RECT 129.650 208.110 129.820 210.510 ;
        RECT 128.070 207.940 129.820 208.110 ;
        RECT 130.170 210.510 131.920 210.680 ;
        RECT 130.170 208.110 130.340 210.510 ;
        RECT 130.880 210.000 131.210 210.170 ;
        RECT 130.740 208.790 130.910 209.830 ;
        RECT 131.180 208.790 131.350 209.830 ;
        RECT 130.880 208.450 131.210 208.620 ;
        RECT 131.750 208.110 131.920 210.510 ;
        RECT 130.170 207.940 131.920 208.110 ;
        RECT 132.280 210.510 137.190 210.680 ;
        RECT 132.280 208.110 132.450 210.510 ;
        RECT 132.990 210.000 133.320 210.170 ;
        RECT 132.850 208.790 133.020 209.830 ;
        RECT 133.290 208.790 133.460 209.830 ;
        RECT 132.990 208.450 133.320 208.620 ;
        RECT 133.860 208.110 134.030 210.510 ;
        RECT 134.570 210.000 134.900 210.170 ;
        RECT 134.430 208.790 134.600 209.830 ;
        RECT 134.870 208.790 135.040 209.830 ;
        RECT 134.570 208.450 134.900 208.620 ;
        RECT 135.440 208.110 135.610 210.510 ;
        RECT 136.150 210.000 136.480 210.170 ;
        RECT 136.010 208.790 136.180 209.830 ;
        RECT 136.450 208.790 136.620 209.830 ;
        RECT 136.150 208.450 136.480 208.620 ;
        RECT 137.020 208.110 137.190 210.510 ;
        RECT 132.280 208.030 137.190 208.110 ;
        RECT 142.820 210.510 144.570 210.680 ;
        RECT 142.820 208.110 142.990 210.510 ;
        RECT 143.530 210.000 143.860 210.170 ;
        RECT 143.390 208.790 143.560 209.830 ;
        RECT 143.830 208.790 144.000 209.830 ;
        RECT 143.530 208.450 143.860 208.620 ;
        RECT 144.400 208.110 144.570 210.510 ;
        RECT 132.280 207.940 137.200 208.030 ;
        RECT 142.820 207.940 144.570 208.110 ;
        RECT 144.920 210.510 146.670 210.680 ;
        RECT 144.920 208.110 145.090 210.510 ;
        RECT 145.630 210.000 145.960 210.170 ;
        RECT 145.490 208.790 145.660 209.830 ;
        RECT 145.930 208.790 146.100 209.830 ;
        RECT 145.630 208.450 145.960 208.620 ;
        RECT 146.500 208.110 146.670 210.510 ;
        RECT 144.920 207.940 146.670 208.110 ;
        RECT 128.090 207.910 129.790 207.940 ;
        RECT 130.190 207.910 131.890 207.940 ;
        RECT 132.360 207.860 137.200 207.940 ;
        RECT 142.840 207.910 144.540 207.940 ;
        RECT 144.940 207.910 146.640 207.940 ;
        RECT 128.090 207.580 129.790 207.610 ;
        RECT 130.190 207.580 131.890 207.610 ;
        RECT 132.360 207.580 137.200 207.660 ;
        RECT 137.630 207.580 142.470 207.660 ;
        RECT 142.840 207.580 144.540 207.610 ;
        RECT 144.940 207.580 146.640 207.610 ;
        RECT 128.070 207.410 129.820 207.580 ;
        RECT 128.070 205.010 128.240 207.410 ;
        RECT 128.780 206.900 129.110 207.070 ;
        RECT 128.640 205.690 128.810 206.730 ;
        RECT 129.080 205.690 129.250 206.730 ;
        RECT 128.780 205.350 129.110 205.520 ;
        RECT 129.650 205.010 129.820 207.410 ;
        RECT 128.070 204.840 129.820 205.010 ;
        RECT 130.170 207.410 131.920 207.580 ;
        RECT 130.170 205.010 130.340 207.410 ;
        RECT 130.880 206.900 131.210 207.070 ;
        RECT 130.740 205.690 130.910 206.730 ;
        RECT 131.180 205.690 131.350 206.730 ;
        RECT 130.880 205.350 131.210 205.520 ;
        RECT 131.750 205.010 131.920 207.410 ;
        RECT 130.170 204.840 131.920 205.010 ;
        RECT 132.280 207.490 137.200 207.580 ;
        RECT 137.550 207.490 142.470 207.580 ;
        RECT 132.280 207.410 137.190 207.490 ;
        RECT 132.280 205.010 132.450 207.410 ;
        RECT 132.990 206.900 133.320 207.070 ;
        RECT 132.850 205.690 133.020 206.730 ;
        RECT 133.290 205.690 133.460 206.730 ;
        RECT 132.990 205.350 133.320 205.520 ;
        RECT 133.860 205.010 134.030 207.410 ;
        RECT 134.570 206.900 134.900 207.070 ;
        RECT 134.430 205.690 134.600 206.730 ;
        RECT 134.870 205.690 135.040 206.730 ;
        RECT 134.570 205.350 134.900 205.520 ;
        RECT 135.440 205.010 135.610 207.410 ;
        RECT 136.150 206.900 136.480 207.070 ;
        RECT 136.010 205.690 136.180 206.730 ;
        RECT 136.450 205.690 136.620 206.730 ;
        RECT 136.150 205.350 136.480 205.520 ;
        RECT 137.020 205.010 137.190 207.410 ;
        RECT 132.280 204.840 137.190 205.010 ;
        RECT 137.550 207.410 142.460 207.490 ;
        RECT 137.550 205.010 137.720 207.410 ;
        RECT 138.260 206.900 138.590 207.070 ;
        RECT 138.120 205.690 138.290 206.730 ;
        RECT 138.560 205.690 138.730 206.730 ;
        RECT 138.260 205.350 138.590 205.520 ;
        RECT 139.130 205.010 139.300 207.410 ;
        RECT 139.840 206.900 140.170 207.070 ;
        RECT 139.700 205.690 139.870 206.730 ;
        RECT 140.140 205.690 140.310 206.730 ;
        RECT 139.840 205.350 140.170 205.520 ;
        RECT 140.710 205.010 140.880 207.410 ;
        RECT 141.420 206.900 141.750 207.070 ;
        RECT 141.280 205.690 141.450 206.730 ;
        RECT 141.720 205.690 141.890 206.730 ;
        RECT 141.420 205.350 141.750 205.520 ;
        RECT 142.290 205.010 142.460 207.410 ;
        RECT 137.550 204.840 142.460 205.010 ;
        RECT 142.820 207.410 144.570 207.580 ;
        RECT 142.820 205.010 142.990 207.410 ;
        RECT 143.530 206.900 143.860 207.070 ;
        RECT 143.390 205.690 143.560 206.730 ;
        RECT 143.830 205.690 144.000 206.730 ;
        RECT 143.530 205.350 143.860 205.520 ;
        RECT 144.400 205.010 144.570 207.410 ;
        RECT 142.820 204.840 144.570 205.010 ;
        RECT 144.920 207.410 146.670 207.580 ;
        RECT 144.920 205.010 145.090 207.410 ;
        RECT 145.630 206.900 145.960 207.070 ;
        RECT 145.490 205.690 145.660 206.730 ;
        RECT 145.930 205.690 146.100 206.730 ;
        RECT 145.630 205.350 145.960 205.520 ;
        RECT 146.500 205.010 146.670 207.410 ;
        RECT 144.920 204.840 146.670 205.010 ;
        RECT 100.710 203.530 125.970 203.700 ;
        RECT 128.070 204.310 129.820 204.480 ;
        RECT 60.740 201.350 71.930 201.520 ;
        RECT 60.740 194.660 60.910 201.350 ;
        RECT 61.390 195.140 63.550 200.870 ;
        RECT 69.120 195.140 71.280 200.870 ;
        RECT 71.760 194.660 71.930 201.350 ;
        RECT 73.910 201.860 99.160 202.030 ;
        RECT 73.910 200.010 74.080 201.860 ;
        RECT 74.760 201.290 78.800 201.460 ;
        RECT 74.420 200.230 74.590 201.230 ;
        RECT 78.970 200.230 79.140 201.230 ;
        RECT 74.840 200.170 78.720 200.200 ;
        RECT 74.760 200.010 78.800 200.170 ;
        RECT 79.480 200.010 79.650 201.860 ;
        RECT 80.610 201.290 85.650 201.460 ;
        RECT 80.270 200.230 80.440 201.230 ;
        RECT 85.820 200.230 85.990 201.230 ;
        RECT 80.610 200.010 85.650 200.170 ;
        RECT 86.450 200.010 86.620 201.860 ;
        RECT 87.580 201.290 92.620 201.460 ;
        RECT 87.240 200.230 87.410 201.230 ;
        RECT 92.790 200.230 92.960 201.230 ;
        RECT 87.580 200.010 92.620 200.170 ;
        RECT 93.420 200.010 93.590 201.860 ;
        RECT 94.270 201.290 98.310 201.460 ;
        RECT 93.930 200.230 94.100 201.230 ;
        RECT 98.480 200.230 98.650 201.230 ;
        RECT 94.350 200.170 98.230 200.200 ;
        RECT 94.270 200.010 98.310 200.170 ;
        RECT 98.990 200.010 99.160 201.860 ;
        RECT 100.720 201.860 125.970 202.030 ;
        RECT 100.720 200.010 100.890 201.860 ;
        RECT 101.570 201.290 105.610 201.460 ;
        RECT 101.230 200.230 101.400 201.230 ;
        RECT 105.780 200.230 105.950 201.230 ;
        RECT 101.650 200.170 105.530 200.200 ;
        RECT 101.570 200.010 105.610 200.170 ;
        RECT 106.290 200.010 106.460 201.860 ;
        RECT 107.420 201.290 112.460 201.460 ;
        RECT 107.080 200.230 107.250 201.230 ;
        RECT 112.630 200.230 112.800 201.230 ;
        RECT 107.420 200.010 112.460 200.170 ;
        RECT 113.260 200.010 113.430 201.860 ;
        RECT 114.390 201.290 119.430 201.460 ;
        RECT 114.050 200.230 114.220 201.230 ;
        RECT 119.600 200.230 119.770 201.230 ;
        RECT 114.390 200.010 119.430 200.170 ;
        RECT 120.230 200.010 120.400 201.860 ;
        RECT 121.080 201.290 125.120 201.460 ;
        RECT 120.740 200.230 120.910 201.230 ;
        RECT 125.290 200.230 125.460 201.230 ;
        RECT 121.160 200.170 125.040 200.200 ;
        RECT 121.080 200.010 125.120 200.170 ;
        RECT 125.800 200.010 125.970 201.860 ;
        RECT 128.070 200.820 128.240 204.310 ;
        RECT 128.780 203.800 129.110 203.970 ;
        RECT 128.640 201.545 128.810 203.585 ;
        RECT 129.080 201.545 129.250 203.585 ;
        RECT 128.780 201.160 129.110 201.330 ;
        RECT 129.650 200.820 129.820 204.310 ;
        RECT 128.070 200.650 129.820 200.820 ;
        RECT 130.170 204.310 131.920 204.480 ;
        RECT 130.170 200.820 130.340 204.310 ;
        RECT 130.880 203.800 131.210 203.970 ;
        RECT 130.740 201.545 130.910 203.585 ;
        RECT 131.180 201.545 131.350 203.585 ;
        RECT 130.880 201.160 131.210 201.330 ;
        RECT 131.750 200.820 131.920 204.310 ;
        RECT 130.170 200.650 131.920 200.820 ;
        RECT 132.280 204.310 137.190 204.480 ;
        RECT 132.280 200.820 132.450 204.310 ;
        RECT 132.990 203.800 133.320 203.970 ;
        RECT 132.850 201.545 133.020 203.585 ;
        RECT 133.290 201.545 133.460 203.585 ;
        RECT 132.990 201.160 133.320 201.330 ;
        RECT 133.860 200.820 134.030 204.310 ;
        RECT 134.570 203.800 134.900 203.970 ;
        RECT 134.430 201.545 134.600 203.585 ;
        RECT 134.870 201.545 135.040 203.585 ;
        RECT 134.570 201.160 134.900 201.330 ;
        RECT 135.440 200.820 135.610 204.310 ;
        RECT 136.150 203.800 136.480 203.970 ;
        RECT 136.010 201.545 136.180 203.585 ;
        RECT 136.450 201.545 136.620 203.585 ;
        RECT 136.150 201.160 136.480 201.330 ;
        RECT 137.020 200.820 137.190 204.310 ;
        RECT 132.280 200.650 137.190 200.820 ;
        RECT 137.550 204.310 142.460 204.480 ;
        RECT 137.550 200.820 137.720 204.310 ;
        RECT 138.260 203.800 138.590 203.970 ;
        RECT 138.120 201.545 138.290 203.585 ;
        RECT 138.560 201.545 138.730 203.585 ;
        RECT 138.260 201.160 138.590 201.330 ;
        RECT 139.130 200.820 139.300 204.310 ;
        RECT 139.840 203.800 140.170 203.970 ;
        RECT 139.700 201.545 139.870 203.585 ;
        RECT 140.140 201.545 140.310 203.585 ;
        RECT 139.840 201.160 140.170 201.330 ;
        RECT 140.710 200.820 140.880 204.310 ;
        RECT 141.420 203.800 141.750 203.970 ;
        RECT 141.280 201.545 141.450 203.585 ;
        RECT 141.720 201.545 141.890 203.585 ;
        RECT 141.420 201.160 141.750 201.330 ;
        RECT 142.290 200.820 142.460 204.310 ;
        RECT 137.550 200.650 142.460 200.820 ;
        RECT 142.820 204.310 144.570 204.480 ;
        RECT 142.820 200.820 142.990 204.310 ;
        RECT 143.530 203.800 143.860 203.970 ;
        RECT 143.390 201.545 143.560 203.585 ;
        RECT 143.830 201.545 144.000 203.585 ;
        RECT 143.530 201.160 143.860 201.330 ;
        RECT 144.400 200.820 144.570 204.310 ;
        RECT 142.820 200.650 144.570 200.820 ;
        RECT 144.920 204.310 146.670 204.480 ;
        RECT 144.920 200.820 145.090 204.310 ;
        RECT 145.630 203.800 145.960 203.970 ;
        RECT 145.490 201.545 145.660 203.585 ;
        RECT 145.930 201.545 146.100 203.585 ;
        RECT 145.630 201.160 145.960 201.330 ;
        RECT 146.500 200.820 146.670 204.310 ;
        RECT 144.920 200.650 146.670 200.820 ;
        RECT 128.090 200.610 129.790 200.650 ;
        RECT 130.190 200.610 131.890 200.650 ;
        RECT 142.840 200.610 144.540 200.650 ;
        RECT 144.940 200.610 146.640 200.650 ;
        RECT 128.090 200.290 129.790 200.330 ;
        RECT 130.190 200.290 131.890 200.330 ;
        RECT 142.840 200.290 144.540 200.330 ;
        RECT 144.940 200.290 146.640 200.330 ;
        RECT 73.900 199.430 99.160 200.010 ;
        RECT 73.900 197.170 79.650 199.430 ;
        RECT 80.610 198.860 85.650 199.030 ;
        RECT 80.270 197.800 80.440 198.800 ;
        RECT 85.820 197.800 85.990 198.800 ;
        RECT 80.610 197.570 85.650 197.740 ;
        RECT 86.450 197.170 86.620 199.430 ;
        RECT 87.580 198.860 92.620 199.030 ;
        RECT 87.240 197.800 87.410 198.800 ;
        RECT 92.790 197.800 92.960 198.800 ;
        RECT 87.580 197.570 92.620 197.740 ;
        RECT 93.420 197.170 99.160 199.430 ;
        RECT 73.900 197.000 99.160 197.170 ;
        RECT 100.710 199.430 125.970 200.010 ;
        RECT 100.710 197.170 106.460 199.430 ;
        RECT 107.420 198.860 112.460 199.030 ;
        RECT 107.080 197.800 107.250 198.800 ;
        RECT 112.630 197.800 112.800 198.800 ;
        RECT 107.420 197.570 112.460 197.740 ;
        RECT 113.260 197.170 113.430 199.430 ;
        RECT 114.390 198.860 119.430 199.030 ;
        RECT 114.050 197.800 114.220 198.800 ;
        RECT 119.600 197.800 119.770 198.800 ;
        RECT 114.390 197.570 119.430 197.740 ;
        RECT 120.230 197.170 125.970 199.430 ;
        RECT 100.710 197.000 125.970 197.170 ;
        RECT 128.070 200.120 129.820 200.290 ;
        RECT 60.740 194.490 71.930 194.660 ;
        RECT 60.740 187.800 60.910 194.490 ;
        RECT 61.390 188.280 63.550 194.010 ;
        RECT 69.120 188.280 71.280 194.010 ;
        RECT 71.760 187.800 71.930 194.490 ;
        RECT 73.900 196.470 99.160 196.640 ;
        RECT 73.900 194.210 79.650 196.470 ;
        RECT 80.610 195.900 85.650 196.070 ;
        RECT 80.270 194.840 80.440 195.840 ;
        RECT 85.820 194.840 85.990 195.840 ;
        RECT 80.610 194.610 85.650 194.780 ;
        RECT 86.450 194.210 86.620 196.470 ;
        RECT 87.580 195.900 92.620 196.070 ;
        RECT 87.240 194.840 87.410 195.840 ;
        RECT 92.790 194.840 92.960 195.840 ;
        RECT 87.580 194.610 92.620 194.780 ;
        RECT 93.420 194.210 99.160 196.470 ;
        RECT 73.900 193.630 99.160 194.210 ;
        RECT 100.710 196.470 125.970 196.640 ;
        RECT 100.710 194.210 106.460 196.470 ;
        RECT 107.420 195.900 112.460 196.070 ;
        RECT 107.080 194.840 107.250 195.840 ;
        RECT 112.630 194.840 112.800 195.840 ;
        RECT 107.420 194.610 112.460 194.780 ;
        RECT 113.260 194.210 113.430 196.470 ;
        RECT 114.390 195.900 119.430 196.070 ;
        RECT 114.050 194.840 114.220 195.840 ;
        RECT 119.600 194.840 119.770 195.840 ;
        RECT 114.390 194.610 119.430 194.780 ;
        RECT 120.230 194.210 125.970 196.470 ;
        RECT 128.070 196.630 128.240 200.120 ;
        RECT 128.780 199.610 129.110 199.780 ;
        RECT 128.640 197.355 128.810 199.395 ;
        RECT 129.080 197.355 129.250 199.395 ;
        RECT 128.780 196.970 129.110 197.140 ;
        RECT 129.650 196.630 129.820 200.120 ;
        RECT 128.070 196.460 129.820 196.630 ;
        RECT 130.170 200.120 131.920 200.290 ;
        RECT 130.170 196.630 130.340 200.120 ;
        RECT 130.880 199.610 131.210 199.780 ;
        RECT 130.740 197.355 130.910 199.395 ;
        RECT 131.180 197.355 131.350 199.395 ;
        RECT 130.880 196.970 131.210 197.140 ;
        RECT 131.750 196.630 131.920 200.120 ;
        RECT 130.170 196.460 131.920 196.630 ;
        RECT 132.280 200.120 137.190 200.290 ;
        RECT 132.280 196.630 132.450 200.120 ;
        RECT 132.990 199.610 133.320 199.780 ;
        RECT 132.850 197.355 133.020 199.395 ;
        RECT 133.290 197.355 133.460 199.395 ;
        RECT 132.990 196.970 133.320 197.140 ;
        RECT 133.860 196.630 134.030 200.120 ;
        RECT 134.570 199.610 134.900 199.780 ;
        RECT 134.430 197.355 134.600 199.395 ;
        RECT 134.870 197.355 135.040 199.395 ;
        RECT 134.570 196.970 134.900 197.140 ;
        RECT 135.440 196.630 135.610 200.120 ;
        RECT 136.150 199.610 136.480 199.780 ;
        RECT 136.010 197.355 136.180 199.395 ;
        RECT 136.450 197.355 136.620 199.395 ;
        RECT 136.150 196.970 136.480 197.140 ;
        RECT 137.020 196.630 137.190 200.120 ;
        RECT 132.280 196.460 137.190 196.630 ;
        RECT 142.820 200.120 144.570 200.290 ;
        RECT 142.820 196.630 142.990 200.120 ;
        RECT 143.530 199.610 143.860 199.780 ;
        RECT 143.390 197.355 143.560 199.395 ;
        RECT 143.830 197.355 144.000 199.395 ;
        RECT 143.530 196.970 143.860 197.140 ;
        RECT 144.400 196.630 144.570 200.120 ;
        RECT 142.820 196.460 144.570 196.630 ;
        RECT 144.920 200.120 146.670 200.290 ;
        RECT 144.920 196.630 145.090 200.120 ;
        RECT 145.630 199.610 145.960 199.780 ;
        RECT 145.490 197.355 145.660 199.395 ;
        RECT 145.930 197.355 146.100 199.395 ;
        RECT 145.630 196.970 145.960 197.140 ;
        RECT 146.500 196.630 146.670 200.120 ;
        RECT 144.920 196.460 146.670 196.630 ;
        RECT 100.710 193.630 125.970 194.210 ;
        RECT 73.910 191.780 74.080 193.630 ;
        RECT 74.760 193.470 78.800 193.630 ;
        RECT 74.840 193.440 78.720 193.470 ;
        RECT 74.420 192.410 74.590 193.410 ;
        RECT 78.970 192.410 79.140 193.410 ;
        RECT 74.760 192.180 78.800 192.350 ;
        RECT 79.480 191.780 79.650 193.630 ;
        RECT 80.610 193.470 85.650 193.630 ;
        RECT 80.270 192.410 80.440 193.410 ;
        RECT 85.820 192.410 85.990 193.410 ;
        RECT 80.610 192.180 85.650 192.350 ;
        RECT 86.450 191.780 86.620 193.630 ;
        RECT 87.580 193.470 92.620 193.630 ;
        RECT 87.240 192.410 87.410 193.410 ;
        RECT 92.790 192.410 92.960 193.410 ;
        RECT 87.580 192.180 92.620 192.350 ;
        RECT 93.420 191.780 93.590 193.630 ;
        RECT 94.270 193.470 98.310 193.630 ;
        RECT 94.350 193.440 98.230 193.470 ;
        RECT 93.930 192.410 94.100 193.410 ;
        RECT 98.480 192.410 98.650 193.410 ;
        RECT 94.270 192.180 98.310 192.350 ;
        RECT 98.990 191.780 99.160 193.630 ;
        RECT 73.910 191.610 99.160 191.780 ;
        RECT 100.720 191.780 100.890 193.630 ;
        RECT 101.570 193.470 105.610 193.630 ;
        RECT 101.650 193.440 105.530 193.470 ;
        RECT 101.230 192.410 101.400 193.410 ;
        RECT 105.780 192.410 105.950 193.410 ;
        RECT 101.570 192.180 105.610 192.350 ;
        RECT 106.290 191.780 106.460 193.630 ;
        RECT 107.420 193.470 112.460 193.630 ;
        RECT 107.080 192.410 107.250 193.410 ;
        RECT 112.630 192.410 112.800 193.410 ;
        RECT 107.420 192.180 112.460 192.350 ;
        RECT 113.260 191.780 113.430 193.630 ;
        RECT 114.390 193.470 119.430 193.630 ;
        RECT 114.050 192.410 114.220 193.410 ;
        RECT 119.600 192.410 119.770 193.410 ;
        RECT 114.390 192.180 119.430 192.350 ;
        RECT 120.230 191.780 120.400 193.630 ;
        RECT 121.080 193.470 125.120 193.630 ;
        RECT 121.160 193.440 125.040 193.470 ;
        RECT 120.740 192.410 120.910 193.410 ;
        RECT 125.290 192.410 125.460 193.410 ;
        RECT 121.080 192.180 125.120 192.350 ;
        RECT 125.800 191.780 125.970 193.630 ;
        RECT 128.070 195.930 129.820 196.100 ;
        RECT 128.070 193.530 128.240 195.930 ;
        RECT 128.780 195.420 129.110 195.590 ;
        RECT 128.640 194.210 128.810 195.250 ;
        RECT 129.080 194.210 129.250 195.250 ;
        RECT 128.780 193.870 129.110 194.040 ;
        RECT 129.650 193.530 129.820 195.930 ;
        RECT 128.070 193.360 129.820 193.530 ;
        RECT 130.170 195.930 131.920 196.100 ;
        RECT 130.170 193.530 130.340 195.930 ;
        RECT 130.880 195.420 131.210 195.590 ;
        RECT 130.740 194.210 130.910 195.250 ;
        RECT 131.180 194.210 131.350 195.250 ;
        RECT 130.880 193.870 131.210 194.040 ;
        RECT 131.750 193.530 131.920 195.930 ;
        RECT 130.170 193.360 131.920 193.530 ;
        RECT 132.280 195.930 137.190 196.100 ;
        RECT 132.280 193.530 132.450 195.930 ;
        RECT 132.990 195.420 133.320 195.590 ;
        RECT 132.850 194.210 133.020 195.250 ;
        RECT 133.290 194.210 133.460 195.250 ;
        RECT 132.990 193.870 133.320 194.040 ;
        RECT 133.860 193.530 134.030 195.930 ;
        RECT 134.570 195.420 134.900 195.590 ;
        RECT 134.430 194.210 134.600 195.250 ;
        RECT 134.870 194.210 135.040 195.250 ;
        RECT 134.570 193.870 134.900 194.040 ;
        RECT 135.440 193.530 135.610 195.930 ;
        RECT 136.150 195.420 136.480 195.590 ;
        RECT 136.010 194.210 136.180 195.250 ;
        RECT 136.450 194.210 136.620 195.250 ;
        RECT 136.150 193.870 136.480 194.040 ;
        RECT 137.020 193.530 137.190 195.930 ;
        RECT 132.280 193.450 137.190 193.530 ;
        RECT 142.820 195.930 144.570 196.100 ;
        RECT 142.820 193.530 142.990 195.930 ;
        RECT 143.530 195.420 143.860 195.590 ;
        RECT 143.390 194.210 143.560 195.250 ;
        RECT 143.830 194.210 144.000 195.250 ;
        RECT 143.530 193.870 143.860 194.040 ;
        RECT 144.400 193.530 144.570 195.930 ;
        RECT 132.280 193.360 137.200 193.450 ;
        RECT 142.820 193.360 144.570 193.530 ;
        RECT 144.920 195.930 146.670 196.100 ;
        RECT 144.920 193.530 145.090 195.930 ;
        RECT 145.630 195.420 145.960 195.590 ;
        RECT 145.490 194.210 145.660 195.250 ;
        RECT 145.930 194.210 146.100 195.250 ;
        RECT 145.630 193.870 145.960 194.040 ;
        RECT 146.500 193.530 146.670 195.930 ;
        RECT 144.920 193.360 146.670 193.530 ;
        RECT 128.090 193.330 129.790 193.360 ;
        RECT 130.190 193.330 131.890 193.360 ;
        RECT 132.360 193.280 137.200 193.360 ;
        RECT 142.840 193.330 144.540 193.360 ;
        RECT 144.940 193.330 146.640 193.360 ;
        RECT 128.090 193.000 129.790 193.030 ;
        RECT 130.190 193.000 131.890 193.030 ;
        RECT 100.720 191.610 125.970 191.780 ;
        RECT 128.070 192.830 129.820 193.000 ;
        RECT 128.070 190.430 128.240 192.830 ;
        RECT 128.780 192.320 129.110 192.490 ;
        RECT 128.640 191.110 128.810 192.150 ;
        RECT 129.080 191.110 129.250 192.150 ;
        RECT 128.780 190.770 129.110 190.940 ;
        RECT 129.650 190.430 129.820 192.830 ;
        RECT 128.070 190.260 129.820 190.430 ;
        RECT 130.170 192.830 131.920 193.000 ;
        RECT 130.170 190.430 130.340 192.830 ;
        RECT 130.880 192.320 131.210 192.490 ;
        RECT 130.740 191.110 130.910 192.150 ;
        RECT 131.180 191.110 131.350 192.150 ;
        RECT 130.880 190.770 131.210 190.940 ;
        RECT 131.750 190.430 131.920 192.830 ;
        RECT 130.170 190.260 131.920 190.430 ;
        RECT 60.740 187.630 71.930 187.800 ;
        RECT 60.740 180.940 60.910 187.630 ;
        RECT 61.390 181.420 63.550 187.150 ;
        RECT 69.120 181.420 71.280 187.150 ;
        RECT 71.760 180.940 71.930 187.630 ;
        RECT 60.740 180.770 71.930 180.940 ;
        RECT 60.740 174.080 60.910 180.770 ;
        RECT 61.390 174.560 63.550 180.290 ;
        RECT 69.120 174.560 71.280 180.290 ;
        RECT 71.760 174.080 71.930 180.770 ;
        RECT 73.900 189.940 99.160 190.110 ;
        RECT 73.900 184.870 75.260 189.940 ;
        RECT 75.835 189.440 85.870 189.610 ;
        RECT 75.450 189.030 75.620 189.380 ;
        RECT 86.085 189.030 86.255 189.380 ;
        RECT 75.835 188.800 85.870 188.970 ;
        RECT 75.835 188.240 85.870 188.410 ;
        RECT 75.450 187.830 75.620 188.180 ;
        RECT 86.085 187.830 86.255 188.180 ;
        RECT 75.835 187.600 85.870 187.770 ;
        RECT 75.835 187.040 85.870 187.210 ;
        RECT 75.450 186.630 75.620 186.980 ;
        RECT 86.085 186.630 86.255 186.980 ;
        RECT 75.835 186.400 85.870 186.570 ;
        RECT 75.835 185.840 85.870 186.010 ;
        RECT 75.450 185.430 75.620 185.780 ;
        RECT 86.085 185.430 86.255 185.780 ;
        RECT 75.835 185.200 85.870 185.370 ;
        RECT 86.450 184.870 86.620 189.940 ;
        RECT 87.195 189.440 97.230 189.610 ;
        RECT 86.810 189.030 86.980 189.380 ;
        RECT 97.445 189.030 97.615 189.380 ;
        RECT 87.195 188.800 97.230 188.970 ;
        RECT 96.470 188.410 97.190 188.500 ;
        RECT 87.195 188.240 97.230 188.410 ;
        RECT 86.810 187.830 86.980 188.180 ;
        RECT 96.470 188.160 97.190 188.240 ;
        RECT 97.445 187.830 97.615 188.180 ;
        RECT 87.195 187.600 97.230 187.770 ;
        RECT 87.195 187.040 97.230 187.210 ;
        RECT 86.810 186.630 86.980 186.980 ;
        RECT 97.445 186.630 97.615 186.980 ;
        RECT 87.195 186.400 97.230 186.570 ;
        RECT 96.470 186.010 97.190 186.100 ;
        RECT 87.195 185.840 97.230 186.010 ;
        RECT 86.810 185.430 86.980 185.780 ;
        RECT 96.470 185.760 97.190 185.840 ;
        RECT 97.445 185.430 97.615 185.780 ;
        RECT 87.195 185.200 97.230 185.370 ;
        RECT 97.805 184.870 99.160 189.940 ;
        RECT 73.900 183.790 99.160 184.870 ;
        RECT 73.900 181.530 80.900 183.790 ;
        RECT 81.625 183.220 91.665 183.390 ;
        RECT 81.240 182.160 81.410 183.160 ;
        RECT 91.880 182.160 92.050 183.160 ;
        RECT 81.625 181.930 91.665 182.100 ;
        RECT 81.705 181.530 91.585 181.930 ;
        RECT 92.380 181.530 99.160 183.790 ;
        RECT 73.900 180.920 99.160 181.530 ;
        RECT 73.900 178.660 76.970 180.920 ;
        RECT 77.685 180.350 85.725 180.520 ;
        RECT 77.300 179.290 77.470 180.290 ;
        RECT 85.940 179.290 86.110 180.290 ;
        RECT 77.685 179.060 85.725 179.230 ;
        RECT 86.450 178.660 86.620 180.920 ;
        RECT 92.380 180.910 99.160 180.920 ;
        RECT 87.345 180.350 95.385 180.520 ;
        RECT 86.960 179.290 87.130 180.290 ;
        RECT 95.600 179.290 95.770 180.290 ;
        RECT 87.345 179.060 95.385 179.230 ;
        RECT 96.110 178.660 99.160 180.910 ;
        RECT 73.900 178.490 99.160 178.660 ;
        RECT 100.710 189.940 125.970 190.110 ;
        RECT 100.710 184.870 102.070 189.940 ;
        RECT 102.645 189.440 112.680 189.610 ;
        RECT 102.260 189.030 102.430 189.380 ;
        RECT 112.895 189.030 113.065 189.380 ;
        RECT 102.645 188.800 112.680 188.970 ;
        RECT 102.645 188.240 112.680 188.410 ;
        RECT 102.260 187.830 102.430 188.180 ;
        RECT 112.895 187.830 113.065 188.180 ;
        RECT 102.645 187.600 112.680 187.770 ;
        RECT 102.645 187.040 112.680 187.210 ;
        RECT 102.260 186.630 102.430 186.980 ;
        RECT 112.895 186.630 113.065 186.980 ;
        RECT 102.645 186.400 112.680 186.570 ;
        RECT 102.645 185.840 112.680 186.010 ;
        RECT 102.260 185.430 102.430 185.780 ;
        RECT 112.895 185.430 113.065 185.780 ;
        RECT 102.645 185.200 112.680 185.370 ;
        RECT 113.260 184.870 113.430 189.940 ;
        RECT 114.005 189.440 124.040 189.610 ;
        RECT 113.620 189.030 113.790 189.380 ;
        RECT 124.255 189.030 124.425 189.380 ;
        RECT 114.005 188.800 124.040 188.970 ;
        RECT 123.280 188.410 124.000 188.500 ;
        RECT 114.005 188.240 124.040 188.410 ;
        RECT 113.620 187.830 113.790 188.180 ;
        RECT 123.280 188.160 124.000 188.240 ;
        RECT 124.255 187.830 124.425 188.180 ;
        RECT 114.005 187.600 124.040 187.770 ;
        RECT 114.005 187.040 124.040 187.210 ;
        RECT 113.620 186.630 113.790 186.980 ;
        RECT 124.255 186.630 124.425 186.980 ;
        RECT 114.005 186.400 124.040 186.570 ;
        RECT 123.280 186.010 124.000 186.100 ;
        RECT 114.005 185.840 124.040 186.010 ;
        RECT 113.620 185.430 113.790 185.780 ;
        RECT 123.280 185.760 124.000 185.840 ;
        RECT 124.255 185.430 124.425 185.780 ;
        RECT 114.005 185.200 124.040 185.370 ;
        RECT 124.615 184.870 125.970 189.940 ;
        RECT 128.070 189.730 129.820 189.900 ;
        RECT 128.070 186.240 128.240 189.730 ;
        RECT 128.780 189.220 129.110 189.390 ;
        RECT 128.640 186.965 128.810 189.005 ;
        RECT 129.080 186.965 129.250 189.005 ;
        RECT 128.780 186.580 129.110 186.750 ;
        RECT 129.650 186.240 129.820 189.730 ;
        RECT 128.070 186.070 129.820 186.240 ;
        RECT 130.170 189.730 131.920 189.900 ;
        RECT 130.170 186.240 130.340 189.730 ;
        RECT 130.880 189.220 131.210 189.390 ;
        RECT 130.740 186.965 130.910 189.005 ;
        RECT 131.180 186.965 131.350 189.005 ;
        RECT 130.880 186.580 131.210 186.750 ;
        RECT 131.750 186.240 131.920 189.730 ;
        RECT 130.170 186.070 131.920 186.240 ;
        RECT 128.090 186.030 129.790 186.070 ;
        RECT 130.190 186.030 131.890 186.070 ;
        RECT 128.090 185.710 129.790 185.750 ;
        RECT 130.190 185.710 131.890 185.750 ;
        RECT 100.710 183.790 125.970 184.870 ;
        RECT 100.710 181.530 107.710 183.790 ;
        RECT 108.435 183.220 118.475 183.390 ;
        RECT 108.050 182.160 108.220 183.160 ;
        RECT 118.690 182.160 118.860 183.160 ;
        RECT 108.435 181.930 118.475 182.100 ;
        RECT 108.515 181.530 118.395 181.930 ;
        RECT 119.190 181.530 125.970 183.790 ;
        RECT 128.070 185.540 129.820 185.710 ;
        RECT 128.070 182.050 128.240 185.540 ;
        RECT 128.780 185.030 129.110 185.200 ;
        RECT 128.640 182.775 128.810 184.815 ;
        RECT 129.080 182.775 129.250 184.815 ;
        RECT 128.780 182.390 129.110 182.560 ;
        RECT 129.650 182.050 129.820 185.540 ;
        RECT 128.070 181.880 129.820 182.050 ;
        RECT 130.170 185.540 131.920 185.710 ;
        RECT 130.170 182.050 130.340 185.540 ;
        RECT 130.880 185.030 131.210 185.200 ;
        RECT 130.740 182.775 130.910 184.815 ;
        RECT 131.180 182.775 131.350 184.815 ;
        RECT 130.880 182.390 131.210 182.560 ;
        RECT 131.750 182.050 131.920 185.540 ;
        RECT 130.170 181.880 131.920 182.050 ;
        RECT 100.710 180.920 125.970 181.530 ;
        RECT 100.710 178.660 103.780 180.920 ;
        RECT 104.495 180.350 112.535 180.520 ;
        RECT 104.110 179.290 104.280 180.290 ;
        RECT 112.750 179.290 112.920 180.290 ;
        RECT 104.495 179.060 112.535 179.230 ;
        RECT 113.260 178.660 113.430 180.920 ;
        RECT 119.190 180.910 125.970 180.920 ;
        RECT 114.155 180.350 122.195 180.520 ;
        RECT 113.770 179.290 113.940 180.290 ;
        RECT 122.410 179.290 122.580 180.290 ;
        RECT 114.155 179.060 122.195 179.230 ;
        RECT 122.920 178.660 125.970 180.910 ;
        RECT 128.070 181.350 129.820 181.520 ;
        RECT 128.070 178.950 128.240 181.350 ;
        RECT 128.780 180.840 129.110 181.010 ;
        RECT 128.640 179.630 128.810 180.670 ;
        RECT 129.080 179.630 129.250 180.670 ;
        RECT 128.780 179.290 129.110 179.460 ;
        RECT 129.650 178.950 129.820 181.350 ;
        RECT 128.070 178.780 129.820 178.950 ;
        RECT 130.170 181.350 131.920 181.520 ;
        RECT 130.170 178.950 130.340 181.350 ;
        RECT 130.880 180.840 131.210 181.010 ;
        RECT 130.740 179.630 130.910 180.670 ;
        RECT 131.180 179.630 131.350 180.670 ;
        RECT 130.880 179.290 131.210 179.460 ;
        RECT 131.750 178.950 131.920 181.350 ;
        RECT 130.170 178.780 131.920 178.950 ;
        RECT 128.090 178.750 129.790 178.780 ;
        RECT 130.190 178.750 131.890 178.780 ;
        RECT 100.710 178.490 125.970 178.660 ;
        RECT 128.090 178.420 129.790 178.450 ;
        RECT 130.190 178.420 131.890 178.450 ;
        RECT 128.070 178.250 129.820 178.420 ;
        RECT 60.740 173.910 71.930 174.080 ;
        RECT 60.740 167.220 60.910 173.910 ;
        RECT 61.390 167.700 63.550 173.430 ;
        RECT 69.120 167.700 71.280 173.430 ;
        RECT 71.760 167.220 71.930 173.910 ;
        RECT 60.740 167.050 71.930 167.220 ;
        RECT 60.740 160.360 60.910 167.050 ;
        RECT 61.390 160.840 63.550 166.570 ;
        RECT 69.120 160.840 71.280 166.570 ;
        RECT 71.760 160.360 71.930 167.050 ;
        RECT 73.900 177.960 99.160 178.130 ;
        RECT 73.900 175.700 76.970 177.960 ;
        RECT 77.685 177.390 85.725 177.560 ;
        RECT 77.300 176.330 77.470 177.330 ;
        RECT 85.940 176.330 86.110 177.330 ;
        RECT 77.685 176.100 85.725 176.270 ;
        RECT 86.450 175.700 86.620 177.960 ;
        RECT 87.345 177.390 95.385 177.560 ;
        RECT 86.960 176.330 87.130 177.330 ;
        RECT 95.600 176.330 95.770 177.330 ;
        RECT 87.345 176.100 95.385 176.270 ;
        RECT 96.110 175.710 99.160 177.960 ;
        RECT 92.380 175.700 99.160 175.710 ;
        RECT 73.900 175.090 99.160 175.700 ;
        RECT 73.900 172.830 80.900 175.090 ;
        RECT 81.705 174.690 91.585 175.090 ;
        RECT 81.625 174.520 91.665 174.690 ;
        RECT 81.240 173.460 81.410 174.460 ;
        RECT 91.880 173.460 92.050 174.460 ;
        RECT 81.625 173.230 91.665 173.400 ;
        RECT 92.380 172.830 99.160 175.090 ;
        RECT 73.900 171.750 99.160 172.830 ;
        RECT 73.900 166.680 75.260 171.750 ;
        RECT 75.835 171.250 85.870 171.420 ;
        RECT 75.450 170.840 75.620 171.190 ;
        RECT 86.085 170.840 86.255 171.190 ;
        RECT 75.835 170.610 85.870 170.780 ;
        RECT 75.835 170.050 85.870 170.220 ;
        RECT 75.450 169.640 75.620 169.990 ;
        RECT 86.085 169.640 86.255 169.990 ;
        RECT 75.835 169.410 85.870 169.580 ;
        RECT 75.835 168.850 85.870 169.020 ;
        RECT 75.450 168.440 75.620 168.790 ;
        RECT 86.085 168.440 86.255 168.790 ;
        RECT 75.835 168.210 85.870 168.380 ;
        RECT 75.835 167.650 85.870 167.820 ;
        RECT 75.450 167.240 75.620 167.590 ;
        RECT 86.085 167.240 86.255 167.590 ;
        RECT 75.835 167.010 85.870 167.180 ;
        RECT 86.450 166.680 86.620 171.750 ;
        RECT 87.195 171.250 97.230 171.420 ;
        RECT 86.810 170.840 86.980 171.190 ;
        RECT 96.470 170.780 97.190 170.860 ;
        RECT 97.445 170.840 97.615 171.190 ;
        RECT 87.195 170.610 97.230 170.780 ;
        RECT 96.470 170.520 97.190 170.610 ;
        RECT 87.195 170.050 97.230 170.220 ;
        RECT 86.810 169.640 86.980 169.990 ;
        RECT 97.445 169.640 97.615 169.990 ;
        RECT 87.195 169.410 97.230 169.580 ;
        RECT 87.195 168.850 97.230 169.020 ;
        RECT 86.810 168.440 86.980 168.790 ;
        RECT 96.470 168.380 97.190 168.460 ;
        RECT 97.445 168.440 97.615 168.790 ;
        RECT 87.195 168.210 97.230 168.380 ;
        RECT 96.470 168.120 97.190 168.210 ;
        RECT 87.195 167.650 97.230 167.820 ;
        RECT 86.810 167.240 86.980 167.590 ;
        RECT 97.445 167.240 97.615 167.590 ;
        RECT 87.195 167.010 97.230 167.180 ;
        RECT 97.805 166.680 99.160 171.750 ;
        RECT 73.900 166.510 99.160 166.680 ;
        RECT 100.710 177.960 125.970 178.130 ;
        RECT 100.710 175.700 103.780 177.960 ;
        RECT 104.495 177.390 112.535 177.560 ;
        RECT 104.110 176.330 104.280 177.330 ;
        RECT 112.750 176.330 112.920 177.330 ;
        RECT 104.495 176.100 112.535 176.270 ;
        RECT 113.260 175.700 113.430 177.960 ;
        RECT 114.155 177.390 122.195 177.560 ;
        RECT 113.770 176.330 113.940 177.330 ;
        RECT 122.410 176.330 122.580 177.330 ;
        RECT 114.155 176.100 122.195 176.270 ;
        RECT 122.920 175.710 125.970 177.960 ;
        RECT 119.190 175.700 125.970 175.710 ;
        RECT 100.710 175.090 125.970 175.700 ;
        RECT 128.070 175.850 128.240 178.250 ;
        RECT 128.780 177.740 129.110 177.910 ;
        RECT 128.640 176.530 128.810 177.570 ;
        RECT 129.080 176.530 129.250 177.570 ;
        RECT 128.780 176.190 129.110 176.360 ;
        RECT 129.650 175.850 129.820 178.250 ;
        RECT 128.070 175.680 129.820 175.850 ;
        RECT 130.170 178.250 131.920 178.420 ;
        RECT 130.170 175.850 130.340 178.250 ;
        RECT 130.880 177.740 131.210 177.910 ;
        RECT 130.740 176.530 130.910 177.570 ;
        RECT 131.180 176.530 131.350 177.570 ;
        RECT 130.880 176.190 131.210 176.360 ;
        RECT 131.750 175.850 131.920 178.250 ;
        RECT 130.170 175.680 131.920 175.850 ;
        RECT 100.710 172.830 107.710 175.090 ;
        RECT 108.515 174.690 118.395 175.090 ;
        RECT 108.435 174.520 118.475 174.690 ;
        RECT 108.050 173.460 108.220 174.460 ;
        RECT 118.690 173.460 118.860 174.460 ;
        RECT 108.435 173.230 118.475 173.400 ;
        RECT 119.190 172.830 125.970 175.090 ;
        RECT 100.710 171.750 125.970 172.830 ;
        RECT 100.710 166.680 102.070 171.750 ;
        RECT 102.645 171.250 112.680 171.420 ;
        RECT 102.260 170.840 102.430 171.190 ;
        RECT 112.895 170.840 113.065 171.190 ;
        RECT 102.645 170.610 112.680 170.780 ;
        RECT 102.645 170.050 112.680 170.220 ;
        RECT 102.260 169.640 102.430 169.990 ;
        RECT 112.895 169.640 113.065 169.990 ;
        RECT 102.645 169.410 112.680 169.580 ;
        RECT 102.645 168.850 112.680 169.020 ;
        RECT 102.260 168.440 102.430 168.790 ;
        RECT 112.895 168.440 113.065 168.790 ;
        RECT 102.645 168.210 112.680 168.380 ;
        RECT 102.645 167.650 112.680 167.820 ;
        RECT 102.260 167.240 102.430 167.590 ;
        RECT 112.895 167.240 113.065 167.590 ;
        RECT 102.645 167.010 112.680 167.180 ;
        RECT 113.260 166.680 113.430 171.750 ;
        RECT 114.005 171.250 124.040 171.420 ;
        RECT 113.620 170.840 113.790 171.190 ;
        RECT 123.280 170.780 124.000 170.860 ;
        RECT 124.255 170.840 124.425 171.190 ;
        RECT 114.005 170.610 124.040 170.780 ;
        RECT 123.280 170.520 124.000 170.610 ;
        RECT 114.005 170.050 124.040 170.220 ;
        RECT 113.620 169.640 113.790 169.990 ;
        RECT 124.255 169.640 124.425 169.990 ;
        RECT 114.005 169.410 124.040 169.580 ;
        RECT 114.005 168.850 124.040 169.020 ;
        RECT 113.620 168.440 113.790 168.790 ;
        RECT 123.280 168.380 124.000 168.460 ;
        RECT 124.255 168.440 124.425 168.790 ;
        RECT 114.005 168.210 124.040 168.380 ;
        RECT 123.280 168.120 124.000 168.210 ;
        RECT 114.005 167.650 124.040 167.820 ;
        RECT 113.620 167.240 113.790 167.590 ;
        RECT 124.255 167.240 124.425 167.590 ;
        RECT 114.005 167.010 124.040 167.180 ;
        RECT 124.615 166.680 125.970 171.750 ;
        RECT 128.070 175.150 129.820 175.320 ;
        RECT 128.070 171.660 128.240 175.150 ;
        RECT 128.780 174.640 129.110 174.810 ;
        RECT 128.640 172.385 128.810 174.425 ;
        RECT 129.080 172.385 129.250 174.425 ;
        RECT 128.780 172.000 129.110 172.170 ;
        RECT 129.650 171.660 129.820 175.150 ;
        RECT 128.070 171.490 129.820 171.660 ;
        RECT 130.170 175.150 131.920 175.320 ;
        RECT 130.170 171.660 130.340 175.150 ;
        RECT 130.880 174.640 131.210 174.810 ;
        RECT 130.740 172.385 130.910 174.425 ;
        RECT 131.180 172.385 131.350 174.425 ;
        RECT 130.880 172.000 131.210 172.170 ;
        RECT 131.750 171.660 131.920 175.150 ;
        RECT 130.170 171.490 131.920 171.660 ;
        RECT 128.090 171.450 129.790 171.490 ;
        RECT 130.190 171.450 131.890 171.490 ;
        RECT 128.090 171.130 129.790 171.170 ;
        RECT 130.190 171.130 131.890 171.170 ;
        RECT 128.070 170.960 129.820 171.130 ;
        RECT 128.070 167.470 128.240 170.960 ;
        RECT 128.780 170.450 129.110 170.620 ;
        RECT 128.640 168.195 128.810 170.235 ;
        RECT 129.080 168.195 129.250 170.235 ;
        RECT 128.780 167.810 129.110 167.980 ;
        RECT 129.650 167.470 129.820 170.960 ;
        RECT 128.070 167.300 129.820 167.470 ;
        RECT 130.170 170.960 131.920 171.130 ;
        RECT 130.170 167.470 130.340 170.960 ;
        RECT 130.880 170.450 131.210 170.620 ;
        RECT 130.740 168.195 130.910 170.235 ;
        RECT 131.180 168.195 131.350 170.235 ;
        RECT 130.880 167.810 131.210 167.980 ;
        RECT 131.750 167.470 131.920 170.960 ;
        RECT 130.170 167.300 131.920 167.470 ;
        RECT 100.710 166.510 125.970 166.680 ;
        RECT 128.070 166.770 129.820 166.940 ;
        RECT 73.910 164.840 99.160 165.010 ;
        RECT 73.910 162.990 74.080 164.840 ;
        RECT 74.760 164.270 78.800 164.440 ;
        RECT 74.420 163.210 74.590 164.210 ;
        RECT 78.970 163.210 79.140 164.210 ;
        RECT 74.840 163.150 78.720 163.180 ;
        RECT 74.760 162.990 78.800 163.150 ;
        RECT 79.480 162.990 79.650 164.840 ;
        RECT 80.610 164.270 85.650 164.440 ;
        RECT 80.270 163.210 80.440 164.210 ;
        RECT 85.820 163.210 85.990 164.210 ;
        RECT 80.610 162.990 85.650 163.150 ;
        RECT 86.450 162.990 86.620 164.840 ;
        RECT 87.580 164.270 92.620 164.440 ;
        RECT 87.240 163.210 87.410 164.210 ;
        RECT 92.790 163.210 92.960 164.210 ;
        RECT 87.580 162.990 92.620 163.150 ;
        RECT 93.420 162.990 93.590 164.840 ;
        RECT 94.270 164.270 98.310 164.440 ;
        RECT 93.930 163.210 94.100 164.210 ;
        RECT 98.480 163.210 98.650 164.210 ;
        RECT 94.350 163.150 98.230 163.180 ;
        RECT 94.270 162.990 98.310 163.150 ;
        RECT 98.990 162.990 99.160 164.840 ;
        RECT 100.720 164.840 125.970 165.010 ;
        RECT 100.720 162.990 100.890 164.840 ;
        RECT 101.570 164.270 105.610 164.440 ;
        RECT 101.230 163.210 101.400 164.210 ;
        RECT 105.780 163.210 105.950 164.210 ;
        RECT 101.650 163.150 105.530 163.180 ;
        RECT 101.570 162.990 105.610 163.150 ;
        RECT 106.290 162.990 106.460 164.840 ;
        RECT 107.420 164.270 112.460 164.440 ;
        RECT 107.080 163.210 107.250 164.210 ;
        RECT 112.630 163.210 112.800 164.210 ;
        RECT 107.420 162.990 112.460 163.150 ;
        RECT 113.260 162.990 113.430 164.840 ;
        RECT 114.390 164.270 119.430 164.440 ;
        RECT 114.050 163.210 114.220 164.210 ;
        RECT 119.600 163.210 119.770 164.210 ;
        RECT 114.390 162.990 119.430 163.150 ;
        RECT 120.230 162.990 120.400 164.840 ;
        RECT 121.080 164.270 125.120 164.440 ;
        RECT 120.740 163.210 120.910 164.210 ;
        RECT 125.290 163.210 125.460 164.210 ;
        RECT 121.160 163.150 125.040 163.180 ;
        RECT 121.080 162.990 125.120 163.150 ;
        RECT 125.800 162.990 125.970 164.840 ;
        RECT 128.070 164.370 128.240 166.770 ;
        RECT 128.780 166.260 129.110 166.430 ;
        RECT 128.640 165.050 128.810 166.090 ;
        RECT 129.080 165.050 129.250 166.090 ;
        RECT 128.780 164.710 129.110 164.880 ;
        RECT 129.650 164.370 129.820 166.770 ;
        RECT 128.070 164.200 129.820 164.370 ;
        RECT 130.170 166.770 131.920 166.940 ;
        RECT 130.170 164.370 130.340 166.770 ;
        RECT 130.880 166.260 131.210 166.430 ;
        RECT 130.740 165.050 130.910 166.090 ;
        RECT 131.180 165.050 131.350 166.090 ;
        RECT 130.880 164.710 131.210 164.880 ;
        RECT 131.750 164.370 131.920 166.770 ;
        RECT 130.170 164.200 131.920 164.370 ;
        RECT 128.090 164.170 129.790 164.200 ;
        RECT 130.190 164.170 131.890 164.200 ;
        RECT 60.740 160.190 71.930 160.360 ;
        RECT 60.740 153.500 60.910 160.190 ;
        RECT 61.390 153.980 63.550 159.710 ;
        RECT 69.120 153.980 71.280 159.710 ;
        RECT 71.760 153.500 71.930 160.190 ;
        RECT 73.900 162.410 99.160 162.990 ;
        RECT 73.900 160.150 79.650 162.410 ;
        RECT 80.610 161.840 85.650 162.010 ;
        RECT 80.270 160.780 80.440 161.780 ;
        RECT 85.820 160.780 85.990 161.780 ;
        RECT 80.610 160.550 85.650 160.720 ;
        RECT 86.450 160.150 86.620 162.410 ;
        RECT 87.580 161.840 92.620 162.010 ;
        RECT 87.240 160.780 87.410 161.780 ;
        RECT 92.790 160.780 92.960 161.780 ;
        RECT 87.580 160.550 92.620 160.720 ;
        RECT 93.420 160.150 99.160 162.410 ;
        RECT 73.900 159.980 99.160 160.150 ;
        RECT 100.710 162.410 125.970 162.990 ;
        RECT 100.710 160.150 106.460 162.410 ;
        RECT 107.420 161.840 112.460 162.010 ;
        RECT 107.080 160.780 107.250 161.780 ;
        RECT 112.630 160.780 112.800 161.780 ;
        RECT 107.420 160.550 112.460 160.720 ;
        RECT 113.260 160.150 113.430 162.410 ;
        RECT 114.390 161.840 119.430 162.010 ;
        RECT 114.050 160.780 114.220 161.780 ;
        RECT 119.600 160.780 119.770 161.780 ;
        RECT 114.390 160.550 119.430 160.720 ;
        RECT 120.230 160.150 125.970 162.410 ;
        RECT 100.710 159.980 125.970 160.150 ;
        RECT 100.700 159.450 125.960 159.620 ;
        RECT 100.700 157.190 106.450 159.450 ;
        RECT 107.410 158.880 112.450 159.050 ;
        RECT 107.070 157.820 107.240 158.820 ;
        RECT 112.620 157.820 112.790 158.820 ;
        RECT 107.410 157.590 112.450 157.760 ;
        RECT 113.250 157.190 113.420 159.450 ;
        RECT 114.380 158.880 119.420 159.050 ;
        RECT 114.040 157.820 114.210 158.820 ;
        RECT 119.590 157.820 119.760 158.820 ;
        RECT 114.380 157.590 119.420 157.760 ;
        RECT 120.220 157.190 125.960 159.450 ;
        RECT 100.700 156.610 125.960 157.190 ;
        RECT 100.710 154.760 100.880 156.610 ;
        RECT 101.560 156.450 105.600 156.610 ;
        RECT 101.640 156.420 105.520 156.450 ;
        RECT 101.220 155.390 101.390 156.390 ;
        RECT 105.770 155.390 105.940 156.390 ;
        RECT 101.560 155.160 105.600 155.330 ;
        RECT 106.280 154.760 106.450 156.610 ;
        RECT 107.410 156.450 112.450 156.610 ;
        RECT 107.070 155.390 107.240 156.390 ;
        RECT 112.620 155.390 112.790 156.390 ;
        RECT 107.410 155.160 112.450 155.330 ;
        RECT 113.250 154.760 113.420 156.610 ;
        RECT 114.380 156.450 119.420 156.610 ;
        RECT 114.040 155.390 114.210 156.390 ;
        RECT 119.590 155.390 119.760 156.390 ;
        RECT 114.380 155.160 119.420 155.330 ;
        RECT 120.220 154.760 120.390 156.610 ;
        RECT 121.070 156.450 125.110 156.610 ;
        RECT 121.150 156.420 125.030 156.450 ;
        RECT 120.730 155.390 120.900 156.390 ;
        RECT 125.280 155.390 125.450 156.390 ;
        RECT 121.070 155.160 125.110 155.330 ;
        RECT 125.790 154.760 125.960 156.610 ;
        RECT 100.710 154.590 125.960 154.760 ;
        RECT 84.190 154.110 86.790 154.230 ;
        RECT 87.060 154.110 97.390 154.230 ;
        RECT 84.190 154.060 97.390 154.110 ;
        RECT 84.190 154.050 84.360 154.060 ;
        RECT 60.740 153.330 71.930 153.500 ;
        RECT 60.740 146.660 60.910 153.330 ;
        RECT 61.390 147.120 63.550 152.850 ;
        RECT 69.120 147.120 71.280 152.850 ;
        RECT 71.760 146.660 71.930 153.330 ;
        RECT 84.150 147.660 84.360 154.050 ;
        RECT 84.990 153.550 85.990 153.720 ;
        RECT 84.760 148.340 84.930 153.380 ;
        RECT 86.050 148.340 86.220 153.380 ;
        RECT 84.990 148.000 85.990 148.170 ;
        RECT 86.620 147.660 87.230 154.060 ;
        RECT 87.710 151.420 89.120 153.580 ;
        RECT 84.150 147.650 87.230 147.660 ;
        RECT 84.150 147.630 86.790 147.650 ;
        RECT 84.190 147.490 86.790 147.630 ;
        RECT 60.740 146.470 71.930 146.660 ;
        RECT 60.750 146.450 71.850 146.470 ;
        RECT 87.060 141.940 87.230 147.650 ;
        RECT 87.710 142.420 89.120 144.580 ;
        RECT 89.600 141.940 89.770 154.060 ;
        RECT 90.250 151.420 91.660 153.580 ;
        RECT 90.250 142.420 91.660 144.580 ;
        RECT 92.140 141.940 92.310 154.060 ;
        RECT 92.790 151.420 94.200 153.580 ;
        RECT 92.790 142.420 94.200 144.580 ;
        RECT 94.680 141.940 94.850 154.060 ;
        RECT 95.330 151.420 96.740 153.580 ;
        RECT 95.330 142.420 96.740 144.580 ;
        RECT 97.220 141.940 97.390 154.060 ;
        RECT 97.750 153.950 100.350 153.970 ;
        RECT 97.750 153.800 100.370 153.950 ;
        RECT 97.750 142.310 97.920 153.800 ;
        RECT 98.550 153.290 99.550 153.460 ;
        RECT 98.320 143.035 98.490 153.075 ;
        RECT 99.610 143.035 99.780 153.075 ;
        RECT 98.550 142.650 99.550 142.820 ;
        RECT 100.180 142.310 100.370 153.800 ;
        RECT 97.750 142.300 100.370 142.310 ;
        RECT 100.700 152.920 125.960 153.090 ;
        RECT 100.700 147.850 102.060 152.920 ;
        RECT 102.635 152.420 112.670 152.590 ;
        RECT 102.250 152.010 102.420 152.360 ;
        RECT 112.885 152.010 113.055 152.360 ;
        RECT 102.635 151.780 112.670 151.950 ;
        RECT 102.635 151.220 112.670 151.390 ;
        RECT 102.250 150.810 102.420 151.160 ;
        RECT 112.885 150.810 113.055 151.160 ;
        RECT 102.635 150.580 112.670 150.750 ;
        RECT 102.635 150.020 112.670 150.190 ;
        RECT 102.250 149.610 102.420 149.960 ;
        RECT 112.885 149.610 113.055 149.960 ;
        RECT 102.635 149.380 112.670 149.550 ;
        RECT 102.635 148.820 112.670 148.990 ;
        RECT 102.250 148.410 102.420 148.760 ;
        RECT 112.885 148.410 113.055 148.760 ;
        RECT 102.635 148.180 112.670 148.350 ;
        RECT 113.250 147.850 113.420 152.920 ;
        RECT 113.995 152.420 124.030 152.590 ;
        RECT 113.610 152.010 113.780 152.360 ;
        RECT 124.245 152.010 124.415 152.360 ;
        RECT 113.995 151.780 124.030 151.950 ;
        RECT 123.270 151.390 123.990 151.480 ;
        RECT 113.995 151.220 124.030 151.390 ;
        RECT 113.610 150.810 113.780 151.160 ;
        RECT 123.270 151.140 123.990 151.220 ;
        RECT 124.245 150.810 124.415 151.160 ;
        RECT 113.995 150.580 124.030 150.750 ;
        RECT 113.995 150.020 124.030 150.190 ;
        RECT 113.610 149.610 113.780 149.960 ;
        RECT 124.245 149.610 124.415 149.960 ;
        RECT 113.995 149.380 124.030 149.550 ;
        RECT 123.270 148.990 123.990 149.080 ;
        RECT 113.995 148.820 124.030 148.990 ;
        RECT 113.610 148.410 113.780 148.760 ;
        RECT 123.270 148.740 123.990 148.820 ;
        RECT 124.245 148.410 124.415 148.760 ;
        RECT 113.995 148.180 124.030 148.350 ;
        RECT 124.605 147.850 125.960 152.920 ;
        RECT 100.700 146.770 125.960 147.850 ;
        RECT 100.700 144.510 107.700 146.770 ;
        RECT 108.425 146.200 118.465 146.370 ;
        RECT 108.040 145.140 108.210 146.140 ;
        RECT 118.680 145.140 118.850 146.140 ;
        RECT 108.425 144.910 118.465 145.080 ;
        RECT 108.505 144.510 118.385 144.910 ;
        RECT 119.180 144.510 125.960 146.770 ;
        RECT 100.700 143.900 125.960 144.510 ;
        RECT 97.750 142.140 100.350 142.300 ;
        RECT 87.060 141.770 97.390 141.940 ;
        RECT 100.700 141.640 103.770 143.900 ;
        RECT 104.485 143.330 112.525 143.500 ;
        RECT 104.100 142.270 104.270 143.270 ;
        RECT 112.740 142.270 112.910 143.270 ;
        RECT 104.485 142.040 112.525 142.210 ;
        RECT 113.250 141.640 113.420 143.900 ;
        RECT 119.180 143.890 125.960 143.900 ;
        RECT 114.145 143.330 122.185 143.500 ;
        RECT 113.760 142.270 113.930 143.270 ;
        RECT 122.400 142.270 122.570 143.270 ;
        RECT 114.145 142.040 122.185 142.210 ;
        RECT 122.910 141.640 125.960 143.890 ;
        RECT 100.700 141.470 125.960 141.640 ;
      LAYER met1 ;
        RECT 60.560 214.970 72.110 215.420 ;
        RECT 61.390 202.000 63.550 214.970 ;
        RECT 73.730 214.950 99.340 215.330 ;
        RECT 61.390 188.280 63.550 200.870 ;
        RECT 69.120 195.140 71.280 214.590 ;
        RECT 73.730 212.720 76.970 214.950 ;
        RECT 77.765 214.610 85.645 214.950 ;
        RECT 87.425 214.610 95.305 214.950 ;
        RECT 77.705 214.380 85.705 214.610 ;
        RECT 87.365 214.380 95.365 214.610 ;
        RECT 77.270 213.990 77.500 214.330 ;
        RECT 85.910 214.270 86.140 214.330 ;
        RECT 86.930 214.270 87.160 214.330 ;
        RECT 85.910 213.990 87.160 214.270 ;
        RECT 95.570 213.990 95.800 214.330 ;
        RECT 77.270 213.730 95.800 213.990 ;
        RECT 77.270 213.340 77.500 213.730 ;
        RECT 85.910 213.430 87.160 213.730 ;
        RECT 85.910 213.340 86.140 213.430 ;
        RECT 86.930 213.370 87.160 213.430 ;
        RECT 95.570 213.370 95.800 213.730 ;
        RECT 77.270 213.080 86.140 213.340 ;
        RECT 87.370 213.320 95.350 213.340 ;
        RECT 87.365 213.090 95.365 213.320 ;
        RECT 87.370 213.080 95.350 213.090 ;
        RECT 96.100 212.720 99.340 214.950 ;
        RECT 73.730 212.360 99.340 212.720 ;
        RECT 100.540 214.950 126.150 215.330 ;
        RECT 100.540 212.720 103.780 214.950 ;
        RECT 104.575 214.610 112.455 214.950 ;
        RECT 114.235 214.610 122.115 214.950 ;
        RECT 104.515 214.380 112.515 214.610 ;
        RECT 114.175 214.380 122.175 214.610 ;
        RECT 104.080 213.990 104.310 214.330 ;
        RECT 112.720 214.270 112.950 214.330 ;
        RECT 113.740 214.270 113.970 214.330 ;
        RECT 112.720 213.990 113.970 214.270 ;
        RECT 122.380 213.990 122.610 214.330 ;
        RECT 104.080 213.730 122.610 213.990 ;
        RECT 104.080 213.340 104.310 213.730 ;
        RECT 112.720 213.430 113.970 213.730 ;
        RECT 112.720 213.340 112.950 213.430 ;
        RECT 113.740 213.370 113.970 213.430 ;
        RECT 122.380 213.370 122.610 213.730 ;
        RECT 104.080 213.080 112.950 213.340 ;
        RECT 114.180 213.320 122.160 213.340 ;
        RECT 114.175 213.090 122.175 213.320 ;
        RECT 114.180 213.080 122.160 213.090 ;
        RECT 122.910 212.720 126.150 214.950 ;
        RECT 127.890 214.650 146.850 215.050 ;
        RECT 100.540 212.360 126.150 212.720 ;
        RECT 128.090 213.860 128.390 214.650 ;
        RECT 128.790 214.160 129.090 214.460 ;
        RECT 128.610 213.860 128.840 213.955 ;
        RECT 128.090 211.960 128.840 213.860 ;
        RECT 128.610 211.955 128.840 211.960 ;
        RECT 129.050 213.860 129.280 213.955 ;
        RECT 130.190 213.860 130.490 214.650 ;
        RECT 130.890 214.160 131.190 214.460 ;
        RECT 130.710 213.860 130.940 213.955 ;
        RECT 129.050 211.960 129.690 213.860 ;
        RECT 130.190 211.960 130.940 213.860 ;
        RECT 129.050 211.955 129.280 211.960 ;
        RECT 81.645 211.510 91.645 211.740 ;
        RECT 108.455 211.510 118.455 211.740 ;
        RECT 81.210 211.400 81.440 211.460 ;
        RECT 91.850 211.400 92.080 211.460 ;
        RECT 108.020 211.400 108.250 211.460 ;
        RECT 118.660 211.400 118.890 211.460 ;
        RECT 81.140 210.560 81.500 211.400 ;
        RECT 91.780 210.560 92.140 211.400 ;
        RECT 107.950 210.560 108.310 211.400 ;
        RECT 118.590 210.560 118.950 211.400 ;
        RECT 128.790 211.060 129.090 211.760 ;
        RECT 127.890 210.660 129.090 211.060 ;
        RECT 81.210 210.500 81.440 210.560 ;
        RECT 91.850 210.500 92.080 210.560 ;
        RECT 108.020 210.500 108.250 210.560 ;
        RECT 118.660 210.500 118.890 210.560 ;
        RECT 81.655 210.450 91.635 210.480 ;
        RECT 108.465 210.450 118.445 210.480 ;
        RECT 81.645 210.220 91.645 210.450 ;
        RECT 108.455 210.220 118.455 210.450 ;
        RECT 128.790 209.960 129.090 210.660 ;
        RECT 129.490 211.060 129.690 211.960 ;
        RECT 130.710 211.955 130.940 211.960 ;
        RECT 131.150 213.860 131.380 213.955 ;
        RECT 132.260 213.900 132.590 214.650 ;
        RECT 132.990 214.160 134.900 214.440 ;
        RECT 136.150 214.170 136.480 214.440 ;
        RECT 136.170 214.160 136.460 214.170 ;
        RECT 132.820 213.900 133.050 213.955 ;
        RECT 131.150 211.960 131.790 213.860 ;
        RECT 132.260 212.010 133.050 213.900 ;
        RECT 131.150 211.955 131.380 211.960 ;
        RECT 130.890 211.060 131.190 211.760 ;
        RECT 129.490 210.660 131.190 211.060 ;
        RECT 128.610 209.760 128.840 209.810 ;
        RECT 73.730 209.120 98.030 209.380 ;
        RECT 100.540 209.120 124.840 209.380 ;
        RECT 85.140 208.470 85.860 208.510 ;
        RECT 87.220 208.470 87.920 208.480 ;
        RECT 75.855 208.240 85.860 208.470 ;
        RECT 87.215 208.240 97.210 208.470 ;
        RECT 85.140 208.190 85.860 208.240 ;
        RECT 87.220 208.210 88.310 208.240 ;
        RECT 75.400 208.130 75.680 208.190 ;
        RECT 75.050 207.940 75.680 208.130 ;
        RECT 75.050 205.730 75.240 207.940 ;
        RECT 75.400 207.880 75.680 207.940 ;
        RECT 86.040 207.880 86.310 208.190 ;
        RECT 86.760 207.880 87.040 208.190 ;
        RECT 97.400 208.130 97.670 208.190 ;
        RECT 97.840 208.130 98.030 209.120 ;
        RECT 111.950 208.470 112.670 208.510 ;
        RECT 114.030 208.470 114.730 208.480 ;
        RECT 102.665 208.240 112.670 208.470 ;
        RECT 114.025 208.240 124.020 208.470 ;
        RECT 111.950 208.190 112.670 208.240 ;
        RECT 114.030 208.210 115.120 208.240 ;
        RECT 102.210 208.130 102.490 208.190 ;
        RECT 97.400 207.940 98.030 208.130 ;
        RECT 97.400 207.880 97.670 207.940 ;
        RECT 75.880 207.830 76.600 207.870 ;
        RECT 87.210 207.830 88.310 207.840 ;
        RECT 96.470 207.830 97.190 207.880 ;
        RECT 75.855 207.600 85.850 207.830 ;
        RECT 87.210 207.600 97.210 207.830 ;
        RECT 75.880 207.550 76.600 207.600 ;
        RECT 87.210 207.580 88.310 207.600 ;
        RECT 96.470 207.540 97.190 207.600 ;
        RECT 85.140 207.270 85.860 207.310 ;
        RECT 87.220 207.270 87.940 207.320 ;
        RECT 75.855 207.040 85.860 207.270 ;
        RECT 87.215 207.040 97.210 207.270 ;
        RECT 85.140 206.990 85.860 207.040 ;
        RECT 75.380 206.680 75.700 206.990 ;
        RECT 86.000 206.660 86.340 207.010 ;
        RECT 86.730 206.660 87.070 207.010 ;
        RECT 87.220 206.990 87.940 207.040 ;
        RECT 97.370 206.660 97.700 207.020 ;
        RECT 77.080 206.630 77.800 206.660 ;
        RECT 95.270 206.630 95.990 206.640 ;
        RECT 75.855 206.400 85.850 206.630 ;
        RECT 87.215 206.400 97.210 206.630 ;
        RECT 77.080 206.350 77.800 206.400 ;
        RECT 95.270 206.380 95.990 206.400 ;
        RECT 85.140 206.070 85.860 206.110 ;
        RECT 87.220 206.070 87.940 206.120 ;
        RECT 75.855 205.840 85.860 206.070 ;
        RECT 87.215 205.840 97.210 206.070 ;
        RECT 85.140 205.790 85.860 205.840 ;
        RECT 87.220 205.810 88.270 205.840 ;
        RECT 75.400 205.730 75.680 205.790 ;
        RECT 75.050 205.540 75.680 205.730 ;
        RECT 75.050 203.430 75.240 205.540 ;
        RECT 75.400 205.480 75.680 205.540 ;
        RECT 86.040 205.480 86.310 205.790 ;
        RECT 86.760 205.480 87.040 205.790 ;
        RECT 97.400 205.730 97.670 205.790 ;
        RECT 97.840 205.730 98.030 207.940 ;
        RECT 97.400 205.540 98.030 205.730 ;
        RECT 101.860 207.940 102.490 208.130 ;
        RECT 101.860 205.730 102.050 207.940 ;
        RECT 102.210 207.880 102.490 207.940 ;
        RECT 112.850 207.880 113.120 208.190 ;
        RECT 113.570 207.880 113.850 208.190 ;
        RECT 124.210 208.130 124.480 208.190 ;
        RECT 124.650 208.130 124.840 209.120 ;
        RECT 128.090 208.860 128.840 209.760 ;
        RECT 128.090 208.160 128.390 208.860 ;
        RECT 128.610 208.810 128.840 208.860 ;
        RECT 129.050 209.760 129.280 209.810 ;
        RECT 129.490 209.760 129.690 210.660 ;
        RECT 130.890 209.960 131.190 210.660 ;
        RECT 131.590 211.060 131.790 211.960 ;
        RECT 132.820 211.955 133.050 212.010 ;
        RECT 133.260 213.900 133.490 213.955 ;
        RECT 134.400 213.900 134.630 213.955 ;
        RECT 133.260 212.020 133.900 213.900 ;
        RECT 133.260 211.955 133.490 212.020 ;
        RECT 133.010 211.740 133.300 211.750 ;
        RECT 131.590 210.660 131.990 211.060 ;
        RECT 130.710 209.760 130.940 209.810 ;
        RECT 129.050 208.860 129.690 209.760 ;
        RECT 130.190 208.860 130.940 209.760 ;
        RECT 129.050 208.810 129.280 208.860 ;
        RECT 128.790 208.360 129.090 208.660 ;
        RECT 130.190 208.160 130.490 208.860 ;
        RECT 130.710 208.810 130.940 208.860 ;
        RECT 131.150 209.760 131.380 209.810 ;
        RECT 131.590 209.760 131.790 210.660 ;
        RECT 132.990 209.980 133.320 211.740 ;
        RECT 133.640 211.030 133.900 212.020 ;
        RECT 134.080 212.020 134.630 213.900 ;
        RECT 133.610 210.680 133.940 211.030 ;
        RECT 133.010 209.970 133.300 209.980 ;
        RECT 131.150 208.860 131.790 209.760 ;
        RECT 132.820 209.750 133.050 209.810 ;
        RECT 132.230 208.870 133.050 209.750 ;
        RECT 131.150 208.810 131.380 208.860 ;
        RECT 130.890 208.360 131.190 208.660 ;
        RECT 132.230 208.160 132.520 208.870 ;
        RECT 132.820 208.810 133.050 208.870 ;
        RECT 133.260 209.750 133.490 209.810 ;
        RECT 133.640 209.750 133.900 210.680 ;
        RECT 133.260 208.870 133.900 209.750 ;
        RECT 134.080 209.750 134.260 212.020 ;
        RECT 134.400 211.955 134.630 212.020 ;
        RECT 134.840 213.900 135.070 213.955 ;
        RECT 135.980 213.900 136.210 213.955 ;
        RECT 134.840 212.010 136.210 213.900 ;
        RECT 134.840 211.955 135.070 212.010 ;
        RECT 134.570 211.470 134.900 211.750 ;
        RECT 134.570 209.970 134.900 211.020 ;
        RECT 134.400 209.750 134.630 209.810 ;
        RECT 134.080 208.870 134.630 209.750 ;
        RECT 133.260 208.810 133.490 208.870 ;
        RECT 134.400 208.810 134.630 208.870 ;
        RECT 134.840 209.750 135.070 209.810 ;
        RECT 135.210 209.750 135.840 212.010 ;
        RECT 135.980 211.955 136.210 212.010 ;
        RECT 136.420 213.900 136.650 213.955 ;
        RECT 136.420 212.010 137.070 213.900 ;
        RECT 136.420 211.955 136.650 212.010 ;
        RECT 136.150 210.700 136.480 211.750 ;
        RECT 136.150 209.990 136.480 210.250 ;
        RECT 136.170 209.970 136.460 209.990 ;
        RECT 135.980 209.750 136.210 209.810 ;
        RECT 134.840 208.870 136.210 209.750 ;
        RECT 134.840 208.810 135.070 208.870 ;
        RECT 135.980 208.810 136.210 208.870 ;
        RECT 136.420 209.750 136.650 209.810 ;
        RECT 136.790 209.750 137.070 212.010 ;
        RECT 142.840 213.860 143.140 214.650 ;
        RECT 143.540 214.160 143.840 214.460 ;
        RECT 143.360 213.860 143.590 213.955 ;
        RECT 142.840 211.960 143.590 213.860 ;
        RECT 143.360 211.955 143.590 211.960 ;
        RECT 143.800 213.860 144.030 213.955 ;
        RECT 144.940 213.860 145.240 214.650 ;
        RECT 145.640 214.160 145.940 214.460 ;
        RECT 145.460 213.860 145.690 213.955 ;
        RECT 143.800 211.960 144.440 213.860 ;
        RECT 144.940 211.960 145.690 213.860 ;
        RECT 143.800 211.955 144.030 211.960 ;
        RECT 143.540 211.060 143.840 211.760 ;
        RECT 142.840 210.660 143.840 211.060 ;
        RECT 143.540 209.960 143.840 210.660 ;
        RECT 144.240 211.060 144.440 211.960 ;
        RECT 145.460 211.955 145.690 211.960 ;
        RECT 145.900 213.860 146.130 213.955 ;
        RECT 145.900 211.960 146.540 213.860 ;
        RECT 145.900 211.955 146.130 211.960 ;
        RECT 145.640 211.060 145.940 211.760 ;
        RECT 144.240 210.660 145.940 211.060 ;
        RECT 143.360 209.760 143.590 209.810 ;
        RECT 136.420 208.870 137.070 209.750 ;
        RECT 136.420 208.810 136.650 208.870 ;
        RECT 142.840 208.860 143.590 209.760 ;
        RECT 133.010 208.640 133.300 208.650 ;
        RECT 134.590 208.640 134.880 208.650 ;
        RECT 136.170 208.640 136.460 208.650 ;
        RECT 132.890 208.310 133.420 208.640 ;
        RECT 134.570 208.370 134.900 208.640 ;
        RECT 136.040 208.310 136.570 208.640 ;
        RECT 142.840 208.160 143.140 208.860 ;
        RECT 143.360 208.810 143.590 208.860 ;
        RECT 143.800 209.760 144.030 209.810 ;
        RECT 144.240 209.760 144.440 210.660 ;
        RECT 145.640 209.960 145.940 210.660 ;
        RECT 146.340 211.060 146.540 211.960 ;
        RECT 146.340 210.660 146.800 211.060 ;
        RECT 145.460 209.760 145.690 209.810 ;
        RECT 143.800 208.860 144.440 209.760 ;
        RECT 144.940 208.860 145.690 209.760 ;
        RECT 143.800 208.810 144.030 208.860 ;
        RECT 143.540 208.360 143.840 208.660 ;
        RECT 144.940 208.160 145.240 208.860 ;
        RECT 145.460 208.810 145.690 208.860 ;
        RECT 145.900 209.760 146.130 209.810 ;
        RECT 146.340 209.760 146.540 210.660 ;
        RECT 145.900 208.860 146.540 209.760 ;
        RECT 145.900 208.810 146.130 208.860 ;
        RECT 145.640 208.360 145.940 208.660 ;
        RECT 124.210 207.940 124.840 208.130 ;
        RECT 124.210 207.880 124.480 207.940 ;
        RECT 102.690 207.830 103.410 207.870 ;
        RECT 114.020 207.830 115.120 207.840 ;
        RECT 123.280 207.830 124.000 207.880 ;
        RECT 102.665 207.600 112.660 207.830 ;
        RECT 114.020 207.600 124.020 207.830 ;
        RECT 102.690 207.550 103.410 207.600 ;
        RECT 114.020 207.580 115.120 207.600 ;
        RECT 123.280 207.540 124.000 207.600 ;
        RECT 111.950 207.270 112.670 207.310 ;
        RECT 114.030 207.270 114.750 207.320 ;
        RECT 102.665 207.040 112.670 207.270 ;
        RECT 114.025 207.040 124.020 207.270 ;
        RECT 111.950 206.990 112.670 207.040 ;
        RECT 102.190 206.680 102.510 206.990 ;
        RECT 112.810 206.660 113.150 207.010 ;
        RECT 113.540 206.660 113.880 207.010 ;
        RECT 114.030 206.990 114.750 207.040 ;
        RECT 124.180 206.660 124.510 207.020 ;
        RECT 103.890 206.630 104.610 206.660 ;
        RECT 122.080 206.630 122.800 206.640 ;
        RECT 102.665 206.400 112.660 206.630 ;
        RECT 114.025 206.400 124.020 206.630 ;
        RECT 103.890 206.350 104.610 206.400 ;
        RECT 122.080 206.380 122.800 206.400 ;
        RECT 111.950 206.070 112.670 206.110 ;
        RECT 114.030 206.070 114.750 206.120 ;
        RECT 102.665 205.840 112.670 206.070 ;
        RECT 114.025 205.840 124.020 206.070 ;
        RECT 111.950 205.790 112.670 205.840 ;
        RECT 114.030 205.810 115.080 205.840 ;
        RECT 102.210 205.730 102.490 205.790 ;
        RECT 101.860 205.540 102.490 205.730 ;
        RECT 97.400 205.480 97.670 205.540 ;
        RECT 75.880 205.430 76.600 205.470 ;
        RECT 87.210 205.430 88.270 205.440 ;
        RECT 96.470 205.430 97.190 205.480 ;
        RECT 75.855 205.200 85.850 205.430 ;
        RECT 87.210 205.200 97.210 205.430 ;
        RECT 75.880 205.150 76.600 205.200 ;
        RECT 87.210 205.180 88.270 205.200 ;
        RECT 96.470 205.140 97.190 205.200 ;
        RECT 85.140 204.870 85.860 204.910 ;
        RECT 87.220 204.870 87.940 204.920 ;
        RECT 75.855 204.640 85.860 204.870 ;
        RECT 87.215 204.640 97.210 204.870 ;
        RECT 85.140 204.590 85.860 204.640 ;
        RECT 75.380 204.280 75.700 204.590 ;
        RECT 86.000 204.260 86.340 204.610 ;
        RECT 86.730 204.260 87.070 204.610 ;
        RECT 87.220 204.590 87.940 204.640 ;
        RECT 97.370 204.260 97.700 204.620 ;
        RECT 77.080 204.230 77.800 204.260 ;
        RECT 95.270 204.230 95.990 204.240 ;
        RECT 75.855 204.000 85.850 204.230 ;
        RECT 87.215 204.000 97.210 204.230 ;
        RECT 77.080 203.950 77.800 204.000 ;
        RECT 95.270 203.980 95.990 204.000 ;
        RECT 101.860 203.430 102.050 205.540 ;
        RECT 102.210 205.480 102.490 205.540 ;
        RECT 112.850 205.480 113.120 205.790 ;
        RECT 113.570 205.480 113.850 205.790 ;
        RECT 124.210 205.730 124.480 205.790 ;
        RECT 124.650 205.730 124.840 207.940 ;
        RECT 127.890 207.360 146.850 208.160 ;
        RECT 128.090 206.660 128.390 207.360 ;
        RECT 128.790 206.860 129.090 207.160 ;
        RECT 128.610 206.660 128.840 206.710 ;
        RECT 128.090 205.760 128.840 206.660 ;
        RECT 124.210 205.540 124.840 205.730 ;
        RECT 128.610 205.710 128.840 205.760 ;
        RECT 129.050 206.660 129.280 206.710 ;
        RECT 130.190 206.660 130.490 207.360 ;
        RECT 130.890 206.860 131.190 207.160 ;
        RECT 130.710 206.660 130.940 206.710 ;
        RECT 129.050 205.760 129.690 206.660 ;
        RECT 130.190 205.760 130.940 206.660 ;
        RECT 129.050 205.710 129.280 205.760 ;
        RECT 124.210 205.480 124.480 205.540 ;
        RECT 102.690 205.430 103.410 205.470 ;
        RECT 114.020 205.430 115.080 205.440 ;
        RECT 123.280 205.430 124.000 205.480 ;
        RECT 102.665 205.200 112.660 205.430 ;
        RECT 114.020 205.200 124.020 205.430 ;
        RECT 102.690 205.150 103.410 205.200 ;
        RECT 114.020 205.180 115.080 205.200 ;
        RECT 123.280 205.140 124.000 205.200 ;
        RECT 111.950 204.870 112.670 204.910 ;
        RECT 114.030 204.870 114.750 204.920 ;
        RECT 102.665 204.640 112.670 204.870 ;
        RECT 114.025 204.640 124.020 204.870 ;
        RECT 128.790 204.860 129.090 205.560 ;
        RECT 111.950 204.590 112.670 204.640 ;
        RECT 102.190 204.280 102.510 204.590 ;
        RECT 112.810 204.260 113.150 204.610 ;
        RECT 113.540 204.260 113.880 204.610 ;
        RECT 114.030 204.590 114.750 204.640 ;
        RECT 124.180 204.260 124.510 204.620 ;
        RECT 127.890 204.460 129.090 204.860 ;
        RECT 103.890 204.230 104.610 204.260 ;
        RECT 122.080 204.230 122.800 204.240 ;
        RECT 102.665 204.000 112.660 204.230 ;
        RECT 114.025 204.000 124.020 204.230 ;
        RECT 103.890 203.950 104.610 204.000 ;
        RECT 122.080 203.980 122.800 204.000 ;
        RECT 128.790 203.760 129.090 204.460 ;
        RECT 129.490 204.860 129.690 205.760 ;
        RECT 130.710 205.710 130.940 205.760 ;
        RECT 131.150 206.660 131.380 206.710 ;
        RECT 131.150 205.760 131.790 206.660 ;
        RECT 132.230 206.650 132.520 207.360 ;
        RECT 132.890 206.880 133.420 207.210 ;
        RECT 134.570 206.880 134.900 207.150 ;
        RECT 136.040 206.880 136.570 207.210 ;
        RECT 133.010 206.870 133.300 206.880 ;
        RECT 134.590 206.870 134.880 206.880 ;
        RECT 136.170 206.870 136.460 206.880 ;
        RECT 132.820 206.650 133.050 206.710 ;
        RECT 132.230 205.770 133.050 206.650 ;
        RECT 131.150 205.710 131.380 205.760 ;
        RECT 130.890 204.860 131.190 205.560 ;
        RECT 129.490 204.460 131.190 204.860 ;
        RECT 128.610 203.560 128.840 203.565 ;
        RECT 73.730 203.170 97.700 203.430 ;
        RECT 100.540 203.170 124.510 203.430 ;
        RECT 77.070 202.770 97.190 203.030 ;
        RECT 103.880 202.770 124.000 203.030 ;
        RECT 75.870 202.370 95.990 202.630 ;
        RECT 102.680 202.370 122.800 202.630 ;
        RECT 128.090 201.660 128.840 203.560 ;
        RECT 74.390 201.490 78.770 201.510 ;
        RECT 80.640 201.490 85.620 201.510 ;
        RECT 87.610 201.490 92.590 201.510 ;
        RECT 74.390 201.250 79.170 201.490 ;
        RECT 80.630 201.260 85.630 201.490 ;
        RECT 87.600 201.260 92.600 201.490 ;
        RECT 80.640 201.250 85.620 201.260 ;
        RECT 87.610 201.250 92.590 201.260 ;
        RECT 93.930 201.250 98.680 201.510 ;
        RECT 74.390 200.860 74.620 201.250 ;
        RECT 78.940 201.150 79.170 201.250 ;
        RECT 93.930 201.230 94.290 201.250 ;
        RECT 93.930 201.210 94.130 201.230 ;
        RECT 80.240 201.150 80.470 201.210 ;
        RECT 85.790 201.150 86.020 201.210 ;
        RECT 87.210 201.150 87.440 201.210 ;
        RECT 92.760 201.150 92.990 201.210 ;
        RECT 93.900 201.150 94.130 201.210 ;
        RECT 78.940 200.860 80.470 201.150 ;
        RECT 85.720 200.860 86.080 201.150 ;
        RECT 74.390 200.600 86.080 200.860 ;
        RECT 74.390 200.250 74.620 200.600 ;
        RECT 78.940 200.310 80.470 200.600 ;
        RECT 85.720 200.310 86.080 200.600 ;
        RECT 87.150 200.860 87.510 201.150 ;
        RECT 92.760 200.860 94.130 201.150 ;
        RECT 98.450 200.860 98.680 201.250 ;
        RECT 87.150 200.600 98.680 200.860 ;
        RECT 87.150 200.310 87.510 200.600 ;
        RECT 92.760 200.310 94.130 200.600 ;
        RECT 78.940 200.250 79.170 200.310 ;
        RECT 80.240 200.250 80.470 200.310 ;
        RECT 85.790 200.250 86.020 200.310 ;
        RECT 87.210 200.250 87.440 200.310 ;
        RECT 92.760 200.250 92.990 200.310 ;
        RECT 93.900 200.250 94.130 200.310 ;
        RECT 98.450 200.250 98.680 200.600 ;
        RECT 101.200 201.490 105.580 201.510 ;
        RECT 107.450 201.490 112.430 201.510 ;
        RECT 114.420 201.490 119.400 201.510 ;
        RECT 101.200 201.250 105.980 201.490 ;
        RECT 107.440 201.260 112.440 201.490 ;
        RECT 114.410 201.260 119.410 201.490 ;
        RECT 107.450 201.250 112.430 201.260 ;
        RECT 114.420 201.250 119.400 201.260 ;
        RECT 120.740 201.250 125.490 201.510 ;
        RECT 101.200 200.860 101.430 201.250 ;
        RECT 105.750 201.150 105.980 201.250 ;
        RECT 120.740 201.230 121.100 201.250 ;
        RECT 120.740 201.210 120.940 201.230 ;
        RECT 107.050 201.150 107.280 201.210 ;
        RECT 112.600 201.150 112.830 201.210 ;
        RECT 114.020 201.150 114.250 201.210 ;
        RECT 119.570 201.150 119.800 201.210 ;
        RECT 120.710 201.150 120.940 201.210 ;
        RECT 105.750 200.860 107.280 201.150 ;
        RECT 112.530 200.860 112.890 201.150 ;
        RECT 101.200 200.600 112.890 200.860 ;
        RECT 101.200 200.250 101.430 200.600 ;
        RECT 105.750 200.310 107.280 200.600 ;
        RECT 112.530 200.310 112.890 200.600 ;
        RECT 113.960 200.860 114.320 201.150 ;
        RECT 119.570 200.860 120.940 201.150 ;
        RECT 125.260 200.860 125.490 201.250 ;
        RECT 128.090 200.870 128.390 201.660 ;
        RECT 128.610 201.565 128.840 201.660 ;
        RECT 129.050 203.560 129.280 203.565 ;
        RECT 129.490 203.560 129.690 204.460 ;
        RECT 130.890 203.760 131.190 204.460 ;
        RECT 131.590 204.860 131.790 205.760 ;
        RECT 132.820 205.710 133.050 205.770 ;
        RECT 133.260 206.650 133.490 206.710 ;
        RECT 134.400 206.650 134.630 206.710 ;
        RECT 133.260 205.770 133.900 206.650 ;
        RECT 133.260 205.710 133.490 205.770 ;
        RECT 133.010 205.540 133.300 205.550 ;
        RECT 131.590 204.460 131.990 204.860 ;
        RECT 130.710 203.560 130.940 203.565 ;
        RECT 129.050 201.660 129.690 203.560 ;
        RECT 130.190 201.660 130.940 203.560 ;
        RECT 129.050 201.565 129.280 201.660 ;
        RECT 128.790 201.060 129.090 201.360 ;
        RECT 130.190 200.870 130.490 201.660 ;
        RECT 130.710 201.565 130.940 201.660 ;
        RECT 131.150 203.560 131.380 203.565 ;
        RECT 131.590 203.560 131.790 204.460 ;
        RECT 132.990 203.780 133.320 205.540 ;
        RECT 133.640 204.840 133.900 205.770 ;
        RECT 134.080 205.770 134.630 206.650 ;
        RECT 133.610 204.490 133.940 204.840 ;
        RECT 133.010 203.770 133.300 203.780 ;
        RECT 131.150 201.660 131.790 203.560 ;
        RECT 132.820 203.510 133.050 203.565 ;
        RECT 131.150 201.565 131.380 201.660 ;
        RECT 132.260 201.620 133.050 203.510 ;
        RECT 130.890 201.060 131.190 201.360 ;
        RECT 132.260 200.870 132.590 201.620 ;
        RECT 132.820 201.565 133.050 201.620 ;
        RECT 133.260 203.500 133.490 203.565 ;
        RECT 133.640 203.500 133.900 204.490 ;
        RECT 133.260 201.620 133.900 203.500 ;
        RECT 134.080 203.500 134.260 205.770 ;
        RECT 134.400 205.710 134.630 205.770 ;
        RECT 134.840 206.650 135.070 206.710 ;
        RECT 135.980 206.650 136.210 206.710 ;
        RECT 134.840 205.770 136.210 206.650 ;
        RECT 134.840 205.710 135.070 205.770 ;
        RECT 134.570 204.500 134.900 205.550 ;
        RECT 134.570 203.770 134.900 204.050 ;
        RECT 134.400 203.500 134.630 203.565 ;
        RECT 134.080 201.620 134.630 203.500 ;
        RECT 133.260 201.565 133.490 201.620 ;
        RECT 134.400 201.565 134.630 201.620 ;
        RECT 134.840 203.510 135.070 203.565 ;
        RECT 135.210 203.510 135.840 205.770 ;
        RECT 135.980 205.710 136.210 205.770 ;
        RECT 136.420 206.650 136.650 206.710 ;
        RECT 137.500 206.650 137.790 207.360 ;
        RECT 138.160 206.880 138.690 207.210 ;
        RECT 139.840 206.880 140.170 207.150 ;
        RECT 141.310 206.880 141.840 207.210 ;
        RECT 138.280 206.870 138.570 206.880 ;
        RECT 139.860 206.870 140.150 206.880 ;
        RECT 141.440 206.870 141.730 206.880 ;
        RECT 138.090 206.650 138.320 206.710 ;
        RECT 136.420 205.770 137.070 206.650 ;
        RECT 137.500 205.770 138.320 206.650 ;
        RECT 136.420 205.710 136.650 205.770 ;
        RECT 136.170 205.530 136.460 205.550 ;
        RECT 136.150 205.270 136.480 205.530 ;
        RECT 136.150 203.770 136.480 204.820 ;
        RECT 135.980 203.510 136.210 203.565 ;
        RECT 134.840 201.620 136.210 203.510 ;
        RECT 134.840 201.565 135.070 201.620 ;
        RECT 135.980 201.565 136.210 201.620 ;
        RECT 136.420 203.510 136.650 203.565 ;
        RECT 136.790 203.510 137.070 205.770 ;
        RECT 138.090 205.710 138.320 205.770 ;
        RECT 138.530 206.650 138.760 206.710 ;
        RECT 139.670 206.650 139.900 206.710 ;
        RECT 138.530 205.770 139.170 206.650 ;
        RECT 138.530 205.710 138.760 205.770 ;
        RECT 138.280 205.540 138.570 205.550 ;
        RECT 138.260 203.780 138.590 205.540 ;
        RECT 138.910 204.840 139.170 205.770 ;
        RECT 139.350 205.770 139.900 206.650 ;
        RECT 138.880 204.490 139.210 204.840 ;
        RECT 138.280 203.770 138.570 203.780 ;
        RECT 138.090 203.510 138.320 203.565 ;
        RECT 136.420 201.620 137.070 203.510 ;
        RECT 137.530 201.620 138.320 203.510 ;
        RECT 136.420 201.565 136.650 201.620 ;
        RECT 132.990 201.080 134.900 201.360 ;
        RECT 136.170 201.350 136.460 201.360 ;
        RECT 136.150 201.080 136.480 201.350 ;
        RECT 137.530 200.870 137.860 201.620 ;
        RECT 138.090 201.565 138.320 201.620 ;
        RECT 138.530 203.500 138.760 203.565 ;
        RECT 138.910 203.500 139.170 204.490 ;
        RECT 138.530 201.620 139.170 203.500 ;
        RECT 139.350 203.500 139.530 205.770 ;
        RECT 139.670 205.710 139.900 205.770 ;
        RECT 140.110 206.650 140.340 206.710 ;
        RECT 141.250 206.650 141.480 206.710 ;
        RECT 140.110 205.770 141.480 206.650 ;
        RECT 140.110 205.710 140.340 205.770 ;
        RECT 139.840 204.500 140.170 205.550 ;
        RECT 139.840 203.770 140.170 204.050 ;
        RECT 139.670 203.500 139.900 203.565 ;
        RECT 139.350 201.620 139.900 203.500 ;
        RECT 138.530 201.565 138.760 201.620 ;
        RECT 139.670 201.565 139.900 201.620 ;
        RECT 140.110 203.510 140.340 203.565 ;
        RECT 140.480 203.510 141.110 205.770 ;
        RECT 141.250 205.710 141.480 205.770 ;
        RECT 141.690 206.650 141.920 206.710 ;
        RECT 142.840 206.660 143.140 207.360 ;
        RECT 143.540 206.860 143.840 207.160 ;
        RECT 143.360 206.660 143.590 206.710 ;
        RECT 141.690 205.770 142.340 206.650 ;
        RECT 141.690 205.710 141.920 205.770 ;
        RECT 141.440 205.530 141.730 205.550 ;
        RECT 141.420 205.270 141.750 205.530 ;
        RECT 141.420 203.770 141.750 204.820 ;
        RECT 141.250 203.510 141.480 203.565 ;
        RECT 140.110 201.620 141.480 203.510 ;
        RECT 140.110 201.565 140.340 201.620 ;
        RECT 141.250 201.565 141.480 201.620 ;
        RECT 141.690 203.510 141.920 203.565 ;
        RECT 142.060 203.510 142.340 205.770 ;
        RECT 142.840 205.760 143.590 206.660 ;
        RECT 143.360 205.710 143.590 205.760 ;
        RECT 143.800 206.660 144.030 206.710 ;
        RECT 144.940 206.660 145.240 207.360 ;
        RECT 145.640 206.860 145.940 207.160 ;
        RECT 145.460 206.660 145.690 206.710 ;
        RECT 143.800 205.760 144.440 206.660 ;
        RECT 144.940 205.760 145.690 206.660 ;
        RECT 143.800 205.710 144.030 205.760 ;
        RECT 143.540 204.860 143.840 205.560 ;
        RECT 142.840 204.460 143.840 204.860 ;
        RECT 143.540 203.760 143.840 204.460 ;
        RECT 144.240 204.860 144.440 205.760 ;
        RECT 145.460 205.710 145.690 205.760 ;
        RECT 145.900 206.660 146.130 206.710 ;
        RECT 145.900 205.760 146.540 206.660 ;
        RECT 145.900 205.710 146.130 205.760 ;
        RECT 145.640 204.860 145.940 205.560 ;
        RECT 144.240 204.460 145.940 204.860 ;
        RECT 143.360 203.560 143.590 203.565 ;
        RECT 141.690 201.620 142.340 203.510 ;
        RECT 142.840 201.660 143.590 203.560 ;
        RECT 141.690 201.565 141.920 201.620 ;
        RECT 138.260 201.080 140.170 201.360 ;
        RECT 141.440 201.350 141.730 201.360 ;
        RECT 141.420 201.080 141.750 201.350 ;
        RECT 142.840 200.870 143.140 201.660 ;
        RECT 143.360 201.565 143.590 201.660 ;
        RECT 143.800 203.560 144.030 203.565 ;
        RECT 144.240 203.560 144.440 204.460 ;
        RECT 145.640 203.760 145.940 204.460 ;
        RECT 146.340 204.860 146.540 205.760 ;
        RECT 146.340 204.460 146.800 204.860 ;
        RECT 145.460 203.560 145.690 203.565 ;
        RECT 143.800 201.660 144.440 203.560 ;
        RECT 144.940 201.660 145.690 203.560 ;
        RECT 143.800 201.565 144.030 201.660 ;
        RECT 143.540 201.060 143.840 201.360 ;
        RECT 144.940 200.870 145.240 201.660 ;
        RECT 145.460 201.565 145.690 201.660 ;
        RECT 145.900 203.560 146.130 203.565 ;
        RECT 146.340 203.560 146.540 204.460 ;
        RECT 145.900 201.660 146.540 203.560 ;
        RECT 145.900 201.565 146.130 201.660 ;
        RECT 145.640 201.060 145.940 201.360 ;
        RECT 113.960 200.600 125.490 200.860 ;
        RECT 113.960 200.310 114.320 200.600 ;
        RECT 119.570 200.310 120.940 200.600 ;
        RECT 105.750 200.250 105.980 200.310 ;
        RECT 107.050 200.250 107.280 200.310 ;
        RECT 112.600 200.250 112.830 200.310 ;
        RECT 114.020 200.250 114.250 200.310 ;
        RECT 119.570 200.250 119.800 200.310 ;
        RECT 120.710 200.250 120.940 200.310 ;
        RECT 125.260 200.250 125.490 200.600 ;
        RECT 74.780 199.970 78.780 200.200 ;
        RECT 80.630 199.970 85.630 200.200 ;
        RECT 87.600 199.970 92.600 200.200 ;
        RECT 94.290 199.970 98.290 200.200 ;
        RECT 101.590 199.970 105.590 200.200 ;
        RECT 107.440 199.970 112.440 200.200 ;
        RECT 114.410 199.970 119.410 200.200 ;
        RECT 121.100 199.970 125.100 200.200 ;
        RECT 127.890 200.070 146.850 200.870 ;
        RECT 75.090 199.600 78.460 199.970 ;
        RECT 81.380 199.600 84.750 199.970 ;
        RECT 88.490 199.600 91.860 199.970 ;
        RECT 101.900 199.600 105.270 199.970 ;
        RECT 108.190 199.600 111.560 199.970 ;
        RECT 115.300 199.600 118.670 199.970 ;
        RECT 73.730 199.430 99.340 199.600 ;
        RECT 73.730 197.200 79.650 199.430 ;
        RECT 80.640 199.060 85.620 199.080 ;
        RECT 87.610 199.060 92.590 199.080 ;
        RECT 80.630 198.830 85.630 199.060 ;
        RECT 87.600 198.830 92.600 199.060 ;
        RECT 80.640 198.820 85.620 198.830 ;
        RECT 87.610 198.820 92.590 198.830 ;
        RECT 80.240 198.440 80.470 198.780 ;
        RECT 85.790 198.720 86.020 198.780 ;
        RECT 87.210 198.720 87.440 198.780 ;
        RECT 85.720 198.440 86.080 198.720 ;
        RECT 80.240 198.180 86.080 198.440 ;
        RECT 80.240 197.820 80.470 198.180 ;
        RECT 85.720 197.880 86.080 198.180 ;
        RECT 87.150 198.440 87.510 198.720 ;
        RECT 92.760 198.440 92.990 198.780 ;
        RECT 87.150 198.180 92.990 198.440 ;
        RECT 87.150 197.880 87.510 198.180 ;
        RECT 85.790 197.820 86.020 197.880 ;
        RECT 87.210 197.820 87.440 197.880 ;
        RECT 92.760 197.820 92.990 198.180 ;
        RECT 80.630 197.540 85.630 197.770 ;
        RECT 87.600 197.540 92.600 197.770 ;
        RECT 80.690 197.200 85.570 197.540 ;
        RECT 87.660 197.200 92.540 197.540 ;
        RECT 93.420 197.200 99.340 199.430 ;
        RECT 73.730 196.440 99.340 197.200 ;
        RECT 73.730 194.210 79.650 196.440 ;
        RECT 80.690 196.100 85.570 196.440 ;
        RECT 87.660 196.100 92.540 196.440 ;
        RECT 80.630 195.870 85.630 196.100 ;
        RECT 87.600 195.870 92.600 196.100 ;
        RECT 80.240 195.460 80.470 195.820 ;
        RECT 85.790 195.760 86.020 195.820 ;
        RECT 87.210 195.760 87.440 195.820 ;
        RECT 85.720 195.460 86.080 195.760 ;
        RECT 80.240 195.200 86.080 195.460 ;
        RECT 80.240 194.860 80.470 195.200 ;
        RECT 85.720 194.920 86.080 195.200 ;
        RECT 87.150 195.460 87.510 195.760 ;
        RECT 92.760 195.460 92.990 195.820 ;
        RECT 87.150 195.200 92.990 195.460 ;
        RECT 87.150 194.920 87.510 195.200 ;
        RECT 85.790 194.860 86.020 194.920 ;
        RECT 87.210 194.860 87.440 194.920 ;
        RECT 92.760 194.860 92.990 195.200 ;
        RECT 80.640 194.810 85.620 194.820 ;
        RECT 87.610 194.810 92.590 194.820 ;
        RECT 80.630 194.580 85.630 194.810 ;
        RECT 87.600 194.580 92.600 194.810 ;
        RECT 80.640 194.560 85.620 194.580 ;
        RECT 87.610 194.560 92.590 194.580 ;
        RECT 93.420 194.210 99.340 196.440 ;
        RECT 73.730 194.040 99.340 194.210 ;
        RECT 100.540 199.430 126.150 199.600 ;
        RECT 100.540 197.200 106.460 199.430 ;
        RECT 107.450 199.060 112.430 199.080 ;
        RECT 114.420 199.060 119.400 199.080 ;
        RECT 107.440 198.830 112.440 199.060 ;
        RECT 114.410 198.830 119.410 199.060 ;
        RECT 107.450 198.820 112.430 198.830 ;
        RECT 114.420 198.820 119.400 198.830 ;
        RECT 107.050 198.440 107.280 198.780 ;
        RECT 112.600 198.720 112.830 198.780 ;
        RECT 114.020 198.720 114.250 198.780 ;
        RECT 112.530 198.440 112.890 198.720 ;
        RECT 107.050 198.180 112.890 198.440 ;
        RECT 107.050 197.820 107.280 198.180 ;
        RECT 112.530 197.880 112.890 198.180 ;
        RECT 113.960 198.440 114.320 198.720 ;
        RECT 119.570 198.440 119.800 198.780 ;
        RECT 113.960 198.180 119.800 198.440 ;
        RECT 113.960 197.880 114.320 198.180 ;
        RECT 112.600 197.820 112.830 197.880 ;
        RECT 114.020 197.820 114.250 197.880 ;
        RECT 119.570 197.820 119.800 198.180 ;
        RECT 107.440 197.540 112.440 197.770 ;
        RECT 114.410 197.540 119.410 197.770 ;
        RECT 107.500 197.200 112.380 197.540 ;
        RECT 114.470 197.200 119.350 197.540 ;
        RECT 120.230 197.200 126.150 199.430 ;
        RECT 128.090 199.280 128.390 200.070 ;
        RECT 128.790 199.580 129.090 199.880 ;
        RECT 128.610 199.280 128.840 199.375 ;
        RECT 128.090 197.380 128.840 199.280 ;
        RECT 128.610 197.375 128.840 197.380 ;
        RECT 129.050 199.280 129.280 199.375 ;
        RECT 130.190 199.280 130.490 200.070 ;
        RECT 130.890 199.580 131.190 199.880 ;
        RECT 130.710 199.280 130.940 199.375 ;
        RECT 129.050 197.380 129.690 199.280 ;
        RECT 130.190 197.380 130.940 199.280 ;
        RECT 129.050 197.375 129.280 197.380 ;
        RECT 100.540 196.440 126.150 197.200 ;
        RECT 128.790 196.480 129.090 197.180 ;
        RECT 100.540 194.210 106.460 196.440 ;
        RECT 107.500 196.100 112.380 196.440 ;
        RECT 114.470 196.100 119.350 196.440 ;
        RECT 107.440 195.870 112.440 196.100 ;
        RECT 114.410 195.870 119.410 196.100 ;
        RECT 107.050 195.460 107.280 195.820 ;
        RECT 112.600 195.760 112.830 195.820 ;
        RECT 114.020 195.760 114.250 195.820 ;
        RECT 112.530 195.460 112.890 195.760 ;
        RECT 107.050 195.200 112.890 195.460 ;
        RECT 107.050 194.860 107.280 195.200 ;
        RECT 112.530 194.920 112.890 195.200 ;
        RECT 113.960 195.460 114.320 195.760 ;
        RECT 119.570 195.460 119.800 195.820 ;
        RECT 113.960 195.200 119.800 195.460 ;
        RECT 113.960 194.920 114.320 195.200 ;
        RECT 112.600 194.860 112.830 194.920 ;
        RECT 114.020 194.860 114.250 194.920 ;
        RECT 119.570 194.860 119.800 195.200 ;
        RECT 107.450 194.810 112.430 194.820 ;
        RECT 114.420 194.810 119.400 194.820 ;
        RECT 107.440 194.580 112.440 194.810 ;
        RECT 114.410 194.580 119.410 194.810 ;
        RECT 107.450 194.560 112.430 194.580 ;
        RECT 114.420 194.560 119.400 194.580 ;
        RECT 120.230 194.210 126.150 196.440 ;
        RECT 127.890 196.080 129.090 196.480 ;
        RECT 128.790 195.380 129.090 196.080 ;
        RECT 129.490 196.480 129.690 197.380 ;
        RECT 130.710 197.375 130.940 197.380 ;
        RECT 131.150 199.280 131.380 199.375 ;
        RECT 132.260 199.320 132.590 200.070 ;
        RECT 132.990 199.580 134.900 199.860 ;
        RECT 136.150 199.590 136.480 199.860 ;
        RECT 136.170 199.580 136.460 199.590 ;
        RECT 132.820 199.320 133.050 199.375 ;
        RECT 131.150 197.380 131.790 199.280 ;
        RECT 132.260 197.430 133.050 199.320 ;
        RECT 131.150 197.375 131.380 197.380 ;
        RECT 130.890 196.480 131.190 197.180 ;
        RECT 129.490 196.080 131.190 196.480 ;
        RECT 128.610 195.180 128.840 195.230 ;
        RECT 100.540 194.040 126.150 194.210 ;
        RECT 128.090 194.280 128.840 195.180 ;
        RECT 61.390 174.560 63.550 187.150 ;
        RECT 69.120 181.420 71.280 194.010 ;
        RECT 75.090 193.670 78.460 194.040 ;
        RECT 81.380 193.670 84.750 194.040 ;
        RECT 88.490 193.670 91.860 194.040 ;
        RECT 101.900 193.670 105.270 194.040 ;
        RECT 108.190 193.670 111.560 194.040 ;
        RECT 115.300 193.670 118.670 194.040 ;
        RECT 74.780 193.440 78.780 193.670 ;
        RECT 80.630 193.440 85.630 193.670 ;
        RECT 87.600 193.440 92.600 193.670 ;
        RECT 94.290 193.440 98.290 193.670 ;
        RECT 101.590 193.440 105.590 193.670 ;
        RECT 107.440 193.440 112.440 193.670 ;
        RECT 114.410 193.440 119.410 193.670 ;
        RECT 121.100 193.440 125.100 193.670 ;
        RECT 128.090 193.580 128.390 194.280 ;
        RECT 128.610 194.230 128.840 194.280 ;
        RECT 129.050 195.180 129.280 195.230 ;
        RECT 129.490 195.180 129.690 196.080 ;
        RECT 130.890 195.380 131.190 196.080 ;
        RECT 131.590 196.480 131.790 197.380 ;
        RECT 132.820 197.375 133.050 197.430 ;
        RECT 133.260 199.320 133.490 199.375 ;
        RECT 134.400 199.320 134.630 199.375 ;
        RECT 133.260 197.440 133.900 199.320 ;
        RECT 133.260 197.375 133.490 197.440 ;
        RECT 133.010 197.160 133.300 197.170 ;
        RECT 131.590 196.080 131.990 196.480 ;
        RECT 130.710 195.180 130.940 195.230 ;
        RECT 129.050 194.280 129.690 195.180 ;
        RECT 130.190 194.280 130.940 195.180 ;
        RECT 129.050 194.230 129.280 194.280 ;
        RECT 128.790 193.780 129.090 194.080 ;
        RECT 130.190 193.580 130.490 194.280 ;
        RECT 130.710 194.230 130.940 194.280 ;
        RECT 131.150 195.180 131.380 195.230 ;
        RECT 131.590 195.180 131.790 196.080 ;
        RECT 132.990 195.400 133.320 197.160 ;
        RECT 133.640 196.450 133.900 197.440 ;
        RECT 134.080 197.440 134.630 199.320 ;
        RECT 133.610 196.100 133.940 196.450 ;
        RECT 133.010 195.390 133.300 195.400 ;
        RECT 131.150 194.280 131.790 195.180 ;
        RECT 132.820 195.170 133.050 195.230 ;
        RECT 132.230 194.290 133.050 195.170 ;
        RECT 131.150 194.230 131.380 194.280 ;
        RECT 130.890 193.780 131.190 194.080 ;
        RECT 132.230 193.580 132.520 194.290 ;
        RECT 132.820 194.230 133.050 194.290 ;
        RECT 133.260 195.170 133.490 195.230 ;
        RECT 133.640 195.170 133.900 196.100 ;
        RECT 133.260 194.290 133.900 195.170 ;
        RECT 134.080 195.170 134.260 197.440 ;
        RECT 134.400 197.375 134.630 197.440 ;
        RECT 134.840 199.320 135.070 199.375 ;
        RECT 135.980 199.320 136.210 199.375 ;
        RECT 134.840 197.430 136.210 199.320 ;
        RECT 134.840 197.375 135.070 197.430 ;
        RECT 134.570 196.890 134.900 197.170 ;
        RECT 134.570 195.390 134.900 196.440 ;
        RECT 134.400 195.170 134.630 195.230 ;
        RECT 134.080 194.290 134.630 195.170 ;
        RECT 133.260 194.230 133.490 194.290 ;
        RECT 134.400 194.230 134.630 194.290 ;
        RECT 134.840 195.170 135.070 195.230 ;
        RECT 135.210 195.170 135.840 197.430 ;
        RECT 135.980 197.375 136.210 197.430 ;
        RECT 136.420 199.320 136.650 199.375 ;
        RECT 136.420 197.430 137.070 199.320 ;
        RECT 136.420 197.375 136.650 197.430 ;
        RECT 136.150 196.120 136.480 197.170 ;
        RECT 136.150 195.410 136.480 195.670 ;
        RECT 136.170 195.390 136.460 195.410 ;
        RECT 135.980 195.170 136.210 195.230 ;
        RECT 134.840 194.290 136.210 195.170 ;
        RECT 134.840 194.230 135.070 194.290 ;
        RECT 135.980 194.230 136.210 194.290 ;
        RECT 136.420 195.170 136.650 195.230 ;
        RECT 136.790 195.170 137.070 197.430 ;
        RECT 142.840 199.280 143.140 200.070 ;
        RECT 143.540 199.580 143.840 199.880 ;
        RECT 143.360 199.280 143.590 199.375 ;
        RECT 142.840 197.380 143.590 199.280 ;
        RECT 143.360 197.375 143.590 197.380 ;
        RECT 143.800 199.280 144.030 199.375 ;
        RECT 144.940 199.280 145.240 200.070 ;
        RECT 145.640 199.580 145.940 199.880 ;
        RECT 145.460 199.280 145.690 199.375 ;
        RECT 143.800 197.380 144.440 199.280 ;
        RECT 144.940 197.380 145.690 199.280 ;
        RECT 143.800 197.375 144.030 197.380 ;
        RECT 141.430 196.480 142.110 196.560 ;
        RECT 143.540 196.480 143.840 197.180 ;
        RECT 141.430 196.080 143.840 196.480 ;
        RECT 141.430 195.620 142.110 196.080 ;
        RECT 143.540 195.380 143.840 196.080 ;
        RECT 144.240 196.480 144.440 197.380 ;
        RECT 145.460 197.375 145.690 197.380 ;
        RECT 145.900 199.280 146.130 199.375 ;
        RECT 145.900 197.380 146.540 199.280 ;
        RECT 145.900 197.375 146.130 197.380 ;
        RECT 145.640 196.480 145.940 197.180 ;
        RECT 144.240 196.080 145.940 196.480 ;
        RECT 143.360 195.180 143.590 195.230 ;
        RECT 136.420 194.290 137.070 195.170 ;
        RECT 136.420 194.230 136.650 194.290 ;
        RECT 142.840 194.280 143.590 195.180 ;
        RECT 133.010 194.060 133.300 194.070 ;
        RECT 134.590 194.060 134.880 194.070 ;
        RECT 136.170 194.060 136.460 194.070 ;
        RECT 132.890 193.730 133.420 194.060 ;
        RECT 134.570 193.790 134.900 194.060 ;
        RECT 136.040 193.730 136.570 194.060 ;
        RECT 142.840 193.580 143.140 194.280 ;
        RECT 143.360 194.230 143.590 194.280 ;
        RECT 143.800 195.180 144.030 195.230 ;
        RECT 144.240 195.180 144.440 196.080 ;
        RECT 145.640 195.380 145.940 196.080 ;
        RECT 146.340 196.480 146.540 197.380 ;
        RECT 146.340 196.080 146.800 196.480 ;
        RECT 145.460 195.180 145.690 195.230 ;
        RECT 143.800 194.280 144.440 195.180 ;
        RECT 144.940 194.280 145.690 195.180 ;
        RECT 143.800 194.230 144.030 194.280 ;
        RECT 143.540 193.780 143.840 194.080 ;
        RECT 144.940 193.580 145.240 194.280 ;
        RECT 145.460 194.230 145.690 194.280 ;
        RECT 145.900 195.180 146.130 195.230 ;
        RECT 146.340 195.180 146.540 196.080 ;
        RECT 145.900 194.280 146.540 195.180 ;
        RECT 145.900 194.230 146.130 194.280 ;
        RECT 145.640 193.780 145.940 194.080 ;
        RECT 74.390 193.040 74.620 193.390 ;
        RECT 78.940 193.330 79.170 193.390 ;
        RECT 80.240 193.330 80.470 193.390 ;
        RECT 85.790 193.330 86.020 193.390 ;
        RECT 87.210 193.330 87.440 193.390 ;
        RECT 92.760 193.330 92.990 193.390 ;
        RECT 93.900 193.330 94.130 193.390 ;
        RECT 78.940 193.040 80.470 193.330 ;
        RECT 85.720 193.040 86.080 193.330 ;
        RECT 74.390 192.780 86.080 193.040 ;
        RECT 74.390 192.390 74.620 192.780 ;
        RECT 78.940 192.490 80.470 192.780 ;
        RECT 85.720 192.490 86.080 192.780 ;
        RECT 87.150 193.040 87.510 193.330 ;
        RECT 92.760 193.040 94.130 193.330 ;
        RECT 98.450 193.040 98.680 193.390 ;
        RECT 87.150 192.780 98.680 193.040 ;
        RECT 87.150 192.490 87.510 192.780 ;
        RECT 92.760 192.490 94.130 192.780 ;
        RECT 78.940 192.390 79.170 192.490 ;
        RECT 80.240 192.430 80.470 192.490 ;
        RECT 85.790 192.430 86.020 192.490 ;
        RECT 87.210 192.430 87.440 192.490 ;
        RECT 92.760 192.430 92.990 192.490 ;
        RECT 93.900 192.430 94.130 192.490 ;
        RECT 93.930 192.410 94.130 192.430 ;
        RECT 93.930 192.390 94.290 192.410 ;
        RECT 98.450 192.390 98.680 192.780 ;
        RECT 74.390 192.150 79.170 192.390 ;
        RECT 80.640 192.380 85.620 192.390 ;
        RECT 87.610 192.380 92.590 192.390 ;
        RECT 80.630 192.150 85.630 192.380 ;
        RECT 87.600 192.150 92.600 192.380 ;
        RECT 74.390 192.130 78.770 192.150 ;
        RECT 80.640 192.130 85.620 192.150 ;
        RECT 87.610 192.130 92.590 192.150 ;
        RECT 93.930 192.130 98.680 192.390 ;
        RECT 101.200 193.040 101.430 193.390 ;
        RECT 105.750 193.330 105.980 193.390 ;
        RECT 107.050 193.330 107.280 193.390 ;
        RECT 112.600 193.330 112.830 193.390 ;
        RECT 114.020 193.330 114.250 193.390 ;
        RECT 119.570 193.330 119.800 193.390 ;
        RECT 120.710 193.330 120.940 193.390 ;
        RECT 105.750 193.040 107.280 193.330 ;
        RECT 112.530 193.040 112.890 193.330 ;
        RECT 101.200 192.780 112.890 193.040 ;
        RECT 101.200 192.390 101.430 192.780 ;
        RECT 105.750 192.490 107.280 192.780 ;
        RECT 112.530 192.490 112.890 192.780 ;
        RECT 113.960 193.040 114.320 193.330 ;
        RECT 119.570 193.040 120.940 193.330 ;
        RECT 125.260 193.040 125.490 193.390 ;
        RECT 113.960 192.780 125.490 193.040 ;
        RECT 127.890 192.780 146.850 193.580 ;
        RECT 113.960 192.490 114.320 192.780 ;
        RECT 119.570 192.490 120.940 192.780 ;
        RECT 105.750 192.390 105.980 192.490 ;
        RECT 107.050 192.430 107.280 192.490 ;
        RECT 112.600 192.430 112.830 192.490 ;
        RECT 114.020 192.430 114.250 192.490 ;
        RECT 119.570 192.430 119.800 192.490 ;
        RECT 120.710 192.430 120.940 192.490 ;
        RECT 120.740 192.410 120.940 192.430 ;
        RECT 120.740 192.390 121.100 192.410 ;
        RECT 125.260 192.390 125.490 192.780 ;
        RECT 101.200 192.150 105.980 192.390 ;
        RECT 107.450 192.380 112.430 192.390 ;
        RECT 114.420 192.380 119.400 192.390 ;
        RECT 107.440 192.150 112.440 192.380 ;
        RECT 114.410 192.150 119.410 192.380 ;
        RECT 101.200 192.130 105.580 192.150 ;
        RECT 107.450 192.130 112.430 192.150 ;
        RECT 114.420 192.130 119.400 192.150 ;
        RECT 120.740 192.130 125.490 192.390 ;
        RECT 128.090 192.080 128.390 192.780 ;
        RECT 128.790 192.280 129.090 192.580 ;
        RECT 128.610 192.080 128.840 192.130 ;
        RECT 75.870 191.010 95.990 191.270 ;
        RECT 102.680 191.010 122.800 191.270 ;
        RECT 128.090 191.180 128.840 192.080 ;
        RECT 128.610 191.130 128.840 191.180 ;
        RECT 129.050 192.080 129.280 192.130 ;
        RECT 130.190 192.080 130.490 192.780 ;
        RECT 130.890 192.280 131.190 192.580 ;
        RECT 130.710 192.080 130.940 192.130 ;
        RECT 129.050 191.180 129.690 192.080 ;
        RECT 130.190 191.180 130.940 192.080 ;
        RECT 129.050 191.130 129.280 191.180 ;
        RECT 77.070 190.610 97.190 190.870 ;
        RECT 103.880 190.610 124.000 190.870 ;
        RECT 73.730 190.210 97.700 190.470 ;
        RECT 100.540 190.210 124.510 190.470 ;
        RECT 128.790 190.280 129.090 190.980 ;
        RECT 75.050 188.100 75.240 190.210 ;
        RECT 77.080 189.640 77.800 189.690 ;
        RECT 95.270 189.640 95.990 189.660 ;
        RECT 75.855 189.410 85.850 189.640 ;
        RECT 87.215 189.410 97.210 189.640 ;
        RECT 77.080 189.380 77.800 189.410 ;
        RECT 95.270 189.400 95.990 189.410 ;
        RECT 75.380 189.050 75.700 189.360 ;
        RECT 85.140 189.000 85.860 189.050 ;
        RECT 86.000 189.030 86.340 189.380 ;
        RECT 86.730 189.030 87.070 189.380 ;
        RECT 87.220 189.000 87.940 189.050 ;
        RECT 97.370 189.020 97.700 189.380 ;
        RECT 75.855 188.770 85.860 189.000 ;
        RECT 87.215 188.770 97.210 189.000 ;
        RECT 85.140 188.730 85.860 188.770 ;
        RECT 87.220 188.720 87.940 188.770 ;
        RECT 75.880 188.440 76.600 188.490 ;
        RECT 87.210 188.440 88.270 188.460 ;
        RECT 96.470 188.440 97.190 188.500 ;
        RECT 75.855 188.210 85.850 188.440 ;
        RECT 87.210 188.210 97.210 188.440 ;
        RECT 75.880 188.170 76.600 188.210 ;
        RECT 87.210 188.200 88.270 188.210 ;
        RECT 96.470 188.160 97.190 188.210 ;
        RECT 75.400 188.100 75.680 188.160 ;
        RECT 75.050 187.910 75.680 188.100 ;
        RECT 75.050 185.700 75.240 187.910 ;
        RECT 75.400 187.850 75.680 187.910 ;
        RECT 86.040 187.850 86.310 188.160 ;
        RECT 86.760 187.850 87.040 188.160 ;
        RECT 97.400 188.100 97.670 188.160 ;
        RECT 101.860 188.100 102.050 190.210 ;
        RECT 127.890 189.880 129.090 190.280 ;
        RECT 103.890 189.640 104.610 189.690 ;
        RECT 122.080 189.640 122.800 189.660 ;
        RECT 102.665 189.410 112.660 189.640 ;
        RECT 114.025 189.410 124.020 189.640 ;
        RECT 103.890 189.380 104.610 189.410 ;
        RECT 122.080 189.400 122.800 189.410 ;
        RECT 102.190 189.050 102.510 189.360 ;
        RECT 111.950 189.000 112.670 189.050 ;
        RECT 112.810 189.030 113.150 189.380 ;
        RECT 113.540 189.030 113.880 189.380 ;
        RECT 114.030 189.000 114.750 189.050 ;
        RECT 124.180 189.020 124.510 189.380 ;
        RECT 128.790 189.180 129.090 189.880 ;
        RECT 129.490 190.280 129.690 191.180 ;
        RECT 130.710 191.130 130.940 191.180 ;
        RECT 131.150 192.080 131.380 192.130 ;
        RECT 131.150 191.180 131.790 192.080 ;
        RECT 132.680 191.575 133.680 192.530 ;
        RECT 131.150 191.130 131.380 191.180 ;
        RECT 130.890 190.280 131.190 190.980 ;
        RECT 129.490 189.880 131.190 190.280 ;
        RECT 102.665 188.770 112.670 189.000 ;
        RECT 114.025 188.770 124.020 189.000 ;
        RECT 128.610 188.980 128.840 188.985 ;
        RECT 111.950 188.730 112.670 188.770 ;
        RECT 114.030 188.720 114.750 188.770 ;
        RECT 102.690 188.440 103.410 188.490 ;
        RECT 114.020 188.440 115.080 188.460 ;
        RECT 123.280 188.440 124.000 188.500 ;
        RECT 102.665 188.210 112.660 188.440 ;
        RECT 114.020 188.210 124.020 188.440 ;
        RECT 102.690 188.170 103.410 188.210 ;
        RECT 114.020 188.200 115.080 188.210 ;
        RECT 123.280 188.160 124.000 188.210 ;
        RECT 102.210 188.100 102.490 188.160 ;
        RECT 97.400 187.910 98.030 188.100 ;
        RECT 97.400 187.850 97.670 187.910 ;
        RECT 85.140 187.800 85.860 187.850 ;
        RECT 87.220 187.800 88.270 187.830 ;
        RECT 75.855 187.570 85.860 187.800 ;
        RECT 87.215 187.570 97.210 187.800 ;
        RECT 85.140 187.530 85.860 187.570 ;
        RECT 87.220 187.520 87.940 187.570 ;
        RECT 77.080 187.240 77.800 187.290 ;
        RECT 95.270 187.240 95.990 187.260 ;
        RECT 75.855 187.010 85.850 187.240 ;
        RECT 87.215 187.010 97.210 187.240 ;
        RECT 77.080 186.980 77.800 187.010 ;
        RECT 95.270 187.000 95.990 187.010 ;
        RECT 75.380 186.650 75.700 186.960 ;
        RECT 85.140 186.600 85.860 186.650 ;
        RECT 86.000 186.630 86.340 186.980 ;
        RECT 86.730 186.630 87.070 186.980 ;
        RECT 87.220 186.600 87.940 186.650 ;
        RECT 97.370 186.620 97.700 186.980 ;
        RECT 75.855 186.370 85.860 186.600 ;
        RECT 87.215 186.370 97.210 186.600 ;
        RECT 85.140 186.330 85.860 186.370 ;
        RECT 87.220 186.320 87.940 186.370 ;
        RECT 75.880 186.040 76.600 186.090 ;
        RECT 87.210 186.040 88.310 186.060 ;
        RECT 96.470 186.040 97.190 186.100 ;
        RECT 75.855 185.810 85.850 186.040 ;
        RECT 87.210 185.810 97.210 186.040 ;
        RECT 75.880 185.770 76.600 185.810 ;
        RECT 87.210 185.800 88.310 185.810 ;
        RECT 96.470 185.760 97.190 185.810 ;
        RECT 75.400 185.700 75.680 185.760 ;
        RECT 75.050 185.510 75.680 185.700 ;
        RECT 75.400 185.450 75.680 185.510 ;
        RECT 86.040 185.450 86.310 185.760 ;
        RECT 86.760 185.450 87.040 185.760 ;
        RECT 97.400 185.700 97.670 185.760 ;
        RECT 97.840 185.700 98.030 187.910 ;
        RECT 97.400 185.510 98.030 185.700 ;
        RECT 101.860 187.910 102.490 188.100 ;
        RECT 101.860 185.700 102.050 187.910 ;
        RECT 102.210 187.850 102.490 187.910 ;
        RECT 112.850 187.850 113.120 188.160 ;
        RECT 113.570 187.850 113.850 188.160 ;
        RECT 124.210 188.100 124.480 188.160 ;
        RECT 124.210 187.910 124.840 188.100 ;
        RECT 124.210 187.850 124.480 187.910 ;
        RECT 111.950 187.800 112.670 187.850 ;
        RECT 114.030 187.800 115.080 187.830 ;
        RECT 102.665 187.570 112.670 187.800 ;
        RECT 114.025 187.570 124.020 187.800 ;
        RECT 111.950 187.530 112.670 187.570 ;
        RECT 114.030 187.520 114.750 187.570 ;
        RECT 103.890 187.240 104.610 187.290 ;
        RECT 122.080 187.240 122.800 187.260 ;
        RECT 102.665 187.010 112.660 187.240 ;
        RECT 114.025 187.010 124.020 187.240 ;
        RECT 103.890 186.980 104.610 187.010 ;
        RECT 122.080 187.000 122.800 187.010 ;
        RECT 102.190 186.650 102.510 186.960 ;
        RECT 111.950 186.600 112.670 186.650 ;
        RECT 112.810 186.630 113.150 186.980 ;
        RECT 113.540 186.630 113.880 186.980 ;
        RECT 114.030 186.600 114.750 186.650 ;
        RECT 124.180 186.620 124.510 186.980 ;
        RECT 102.665 186.370 112.670 186.600 ;
        RECT 114.025 186.370 124.020 186.600 ;
        RECT 111.950 186.330 112.670 186.370 ;
        RECT 114.030 186.320 114.750 186.370 ;
        RECT 102.690 186.040 103.410 186.090 ;
        RECT 114.020 186.040 115.120 186.060 ;
        RECT 123.280 186.040 124.000 186.100 ;
        RECT 102.665 185.810 112.660 186.040 ;
        RECT 114.020 185.810 124.020 186.040 ;
        RECT 102.690 185.770 103.410 185.810 ;
        RECT 114.020 185.800 115.120 185.810 ;
        RECT 123.280 185.760 124.000 185.810 ;
        RECT 102.210 185.700 102.490 185.760 ;
        RECT 101.860 185.510 102.490 185.700 ;
        RECT 97.400 185.450 97.670 185.510 ;
        RECT 85.140 185.400 85.860 185.450 ;
        RECT 87.220 185.400 88.310 185.430 ;
        RECT 75.855 185.170 85.860 185.400 ;
        RECT 87.215 185.170 97.210 185.400 ;
        RECT 85.140 185.130 85.860 185.170 ;
        RECT 87.220 185.160 87.920 185.170 ;
        RECT 97.840 184.520 98.030 185.510 ;
        RECT 102.210 185.450 102.490 185.510 ;
        RECT 112.850 185.450 113.120 185.760 ;
        RECT 113.570 185.450 113.850 185.760 ;
        RECT 124.210 185.700 124.480 185.760 ;
        RECT 124.650 185.700 124.840 187.910 ;
        RECT 128.090 187.080 128.840 188.980 ;
        RECT 128.090 186.290 128.390 187.080 ;
        RECT 128.610 186.985 128.840 187.080 ;
        RECT 129.050 188.980 129.280 188.985 ;
        RECT 129.490 188.980 129.690 189.880 ;
        RECT 130.890 189.180 131.190 189.880 ;
        RECT 131.590 190.280 131.790 191.180 ;
        RECT 132.680 190.280 133.680 190.575 ;
        RECT 131.590 189.880 133.680 190.280 ;
        RECT 130.710 188.980 130.940 188.985 ;
        RECT 129.050 187.080 129.690 188.980 ;
        RECT 130.190 187.080 130.940 188.980 ;
        RECT 129.050 186.985 129.280 187.080 ;
        RECT 128.790 186.480 129.090 186.780 ;
        RECT 130.190 186.290 130.490 187.080 ;
        RECT 130.710 186.985 130.940 187.080 ;
        RECT 131.150 188.980 131.380 188.985 ;
        RECT 131.590 188.980 131.790 189.880 ;
        RECT 131.150 187.080 131.790 188.980 ;
        RECT 131.150 186.985 131.380 187.080 ;
        RECT 130.890 186.480 131.190 186.780 ;
        RECT 124.210 185.510 124.840 185.700 ;
        RECT 124.210 185.450 124.480 185.510 ;
        RECT 111.950 185.400 112.670 185.450 ;
        RECT 114.030 185.400 115.120 185.430 ;
        RECT 102.665 185.170 112.670 185.400 ;
        RECT 114.025 185.170 124.020 185.400 ;
        RECT 111.950 185.130 112.670 185.170 ;
        RECT 114.030 185.160 114.730 185.170 ;
        RECT 124.650 184.520 124.840 185.510 ;
        RECT 127.890 185.490 146.850 186.290 ;
        RECT 73.730 184.260 98.030 184.520 ;
        RECT 100.540 184.260 124.840 184.520 ;
        RECT 128.090 184.700 128.390 185.490 ;
        RECT 128.790 185.000 129.090 185.300 ;
        RECT 128.610 184.700 128.840 184.795 ;
        RECT 81.645 183.190 91.645 183.420 ;
        RECT 108.455 183.190 118.455 183.420 ;
        RECT 81.655 183.160 91.635 183.190 ;
        RECT 108.465 183.160 118.445 183.190 ;
        RECT 81.210 183.080 81.440 183.140 ;
        RECT 91.850 183.080 92.080 183.140 ;
        RECT 108.020 183.080 108.250 183.140 ;
        RECT 118.660 183.080 118.890 183.140 ;
        RECT 81.140 182.240 81.500 183.080 ;
        RECT 91.780 182.240 92.140 183.080 ;
        RECT 107.950 182.240 108.310 183.080 ;
        RECT 118.590 182.240 118.950 183.080 ;
        RECT 128.090 182.800 128.840 184.700 ;
        RECT 128.610 182.795 128.840 182.800 ;
        RECT 129.050 184.700 129.280 184.795 ;
        RECT 130.190 184.700 130.490 185.490 ;
        RECT 130.890 185.000 131.190 185.300 ;
        RECT 130.710 184.700 130.940 184.795 ;
        RECT 129.050 182.800 129.690 184.700 ;
        RECT 130.190 182.800 130.940 184.700 ;
        RECT 129.050 182.795 129.280 182.800 ;
        RECT 81.210 182.180 81.440 182.240 ;
        RECT 91.850 182.180 92.080 182.240 ;
        RECT 108.020 182.180 108.250 182.240 ;
        RECT 118.660 182.180 118.890 182.240 ;
        RECT 81.645 181.900 91.645 182.130 ;
        RECT 108.455 181.900 118.455 182.130 ;
        RECT 128.790 181.900 129.090 182.600 ;
        RECT 127.890 181.500 129.090 181.900 ;
        RECT 73.730 180.920 99.340 181.280 ;
        RECT 61.390 160.840 63.550 173.430 ;
        RECT 69.120 167.700 71.280 180.290 ;
        RECT 73.730 178.690 76.970 180.920 ;
        RECT 77.270 180.300 86.140 180.560 ;
        RECT 87.370 180.550 95.350 180.560 ;
        RECT 87.365 180.320 95.365 180.550 ;
        RECT 87.370 180.300 95.350 180.320 ;
        RECT 77.270 179.910 77.500 180.300 ;
        RECT 85.910 180.210 86.140 180.300 ;
        RECT 86.930 180.210 87.160 180.270 ;
        RECT 85.910 179.910 87.160 180.210 ;
        RECT 95.570 179.910 95.800 180.270 ;
        RECT 77.270 179.650 95.800 179.910 ;
        RECT 77.270 179.310 77.500 179.650 ;
        RECT 85.910 179.370 87.160 179.650 ;
        RECT 85.910 179.310 86.140 179.370 ;
        RECT 86.930 179.310 87.160 179.370 ;
        RECT 95.570 179.310 95.800 179.650 ;
        RECT 77.705 179.030 85.705 179.260 ;
        RECT 87.365 179.030 95.365 179.260 ;
        RECT 77.765 178.690 85.645 179.030 ;
        RECT 87.425 178.690 95.305 179.030 ;
        RECT 96.100 178.690 99.340 180.920 ;
        RECT 73.730 177.930 99.340 178.690 ;
        RECT 73.730 175.700 76.970 177.930 ;
        RECT 77.765 177.590 85.645 177.930 ;
        RECT 87.425 177.590 95.305 177.930 ;
        RECT 77.705 177.360 85.705 177.590 ;
        RECT 87.365 177.360 95.365 177.590 ;
        RECT 77.270 176.970 77.500 177.310 ;
        RECT 85.910 177.250 86.140 177.310 ;
        RECT 86.930 177.250 87.160 177.310 ;
        RECT 85.910 176.970 87.160 177.250 ;
        RECT 95.570 176.970 95.800 177.310 ;
        RECT 77.270 176.710 95.800 176.970 ;
        RECT 77.270 176.320 77.500 176.710 ;
        RECT 85.910 176.410 87.160 176.710 ;
        RECT 85.910 176.320 86.140 176.410 ;
        RECT 86.930 176.350 87.160 176.410 ;
        RECT 95.570 176.350 95.800 176.710 ;
        RECT 77.270 176.060 86.140 176.320 ;
        RECT 87.370 176.300 95.350 176.320 ;
        RECT 87.365 176.070 95.365 176.300 ;
        RECT 87.370 176.060 95.350 176.070 ;
        RECT 96.100 175.700 99.340 177.930 ;
        RECT 73.730 175.340 99.340 175.700 ;
        RECT 100.540 180.920 126.150 181.280 ;
        RECT 100.540 178.690 103.780 180.920 ;
        RECT 104.080 180.300 112.950 180.560 ;
        RECT 114.180 180.550 122.160 180.560 ;
        RECT 114.175 180.320 122.175 180.550 ;
        RECT 114.180 180.300 122.160 180.320 ;
        RECT 104.080 179.910 104.310 180.300 ;
        RECT 112.720 180.210 112.950 180.300 ;
        RECT 113.740 180.210 113.970 180.270 ;
        RECT 112.720 179.910 113.970 180.210 ;
        RECT 122.380 179.910 122.610 180.270 ;
        RECT 104.080 179.650 122.610 179.910 ;
        RECT 104.080 179.310 104.310 179.650 ;
        RECT 112.720 179.370 113.970 179.650 ;
        RECT 112.720 179.310 112.950 179.370 ;
        RECT 113.740 179.310 113.970 179.370 ;
        RECT 122.380 179.310 122.610 179.650 ;
        RECT 104.515 179.030 112.515 179.260 ;
        RECT 114.175 179.030 122.175 179.260 ;
        RECT 104.575 178.690 112.455 179.030 ;
        RECT 114.235 178.690 122.115 179.030 ;
        RECT 122.910 178.690 126.150 180.920 ;
        RECT 128.790 180.800 129.090 181.500 ;
        RECT 129.490 181.900 129.690 182.800 ;
        RECT 130.710 182.795 130.940 182.800 ;
        RECT 131.150 184.700 131.380 184.795 ;
        RECT 131.150 182.800 131.790 184.700 ;
        RECT 131.150 182.795 131.380 182.800 ;
        RECT 130.890 181.900 131.190 182.600 ;
        RECT 129.490 181.500 131.190 181.900 ;
        RECT 128.610 180.600 128.840 180.650 ;
        RECT 128.090 179.700 128.840 180.600 ;
        RECT 128.090 179.000 128.390 179.700 ;
        RECT 128.610 179.650 128.840 179.700 ;
        RECT 129.050 180.600 129.280 180.650 ;
        RECT 129.490 180.600 129.690 181.500 ;
        RECT 130.890 180.800 131.190 181.500 ;
        RECT 131.590 181.900 131.790 182.800 ;
        RECT 131.590 181.500 131.990 181.900 ;
        RECT 130.710 180.600 130.940 180.650 ;
        RECT 129.050 179.700 129.690 180.600 ;
        RECT 130.190 179.700 130.940 180.600 ;
        RECT 129.050 179.650 129.280 179.700 ;
        RECT 128.790 179.200 129.090 179.500 ;
        RECT 130.190 179.000 130.490 179.700 ;
        RECT 130.710 179.650 130.940 179.700 ;
        RECT 131.150 180.600 131.380 180.650 ;
        RECT 131.590 180.600 131.790 181.500 ;
        RECT 131.150 179.700 131.790 180.600 ;
        RECT 131.150 179.650 131.380 179.700 ;
        RECT 130.890 179.200 131.190 179.500 ;
        RECT 100.540 177.930 126.150 178.690 ;
        RECT 127.890 178.200 146.850 179.000 ;
        RECT 100.540 175.700 103.780 177.930 ;
        RECT 104.575 177.590 112.455 177.930 ;
        RECT 114.235 177.590 122.115 177.930 ;
        RECT 104.515 177.360 112.515 177.590 ;
        RECT 114.175 177.360 122.175 177.590 ;
        RECT 104.080 176.970 104.310 177.310 ;
        RECT 112.720 177.250 112.950 177.310 ;
        RECT 113.740 177.250 113.970 177.310 ;
        RECT 112.720 176.970 113.970 177.250 ;
        RECT 122.380 176.970 122.610 177.310 ;
        RECT 104.080 176.710 122.610 176.970 ;
        RECT 104.080 176.320 104.310 176.710 ;
        RECT 112.720 176.410 113.970 176.710 ;
        RECT 112.720 176.320 112.950 176.410 ;
        RECT 113.740 176.350 113.970 176.410 ;
        RECT 122.380 176.350 122.610 176.710 ;
        RECT 104.080 176.060 112.950 176.320 ;
        RECT 114.180 176.300 122.160 176.320 ;
        RECT 114.175 176.070 122.175 176.300 ;
        RECT 114.180 176.060 122.160 176.070 ;
        RECT 122.910 175.700 126.150 177.930 ;
        RECT 128.090 177.500 128.390 178.200 ;
        RECT 128.790 177.700 129.090 178.000 ;
        RECT 128.610 177.500 128.840 177.550 ;
        RECT 128.090 176.600 128.840 177.500 ;
        RECT 128.610 176.550 128.840 176.600 ;
        RECT 129.050 177.500 129.280 177.550 ;
        RECT 130.190 177.500 130.490 178.200 ;
        RECT 130.890 177.700 131.190 178.000 ;
        RECT 130.710 177.500 130.940 177.550 ;
        RECT 129.050 176.600 129.690 177.500 ;
        RECT 130.190 176.600 130.940 177.500 ;
        RECT 129.050 176.550 129.280 176.600 ;
        RECT 128.790 175.700 129.090 176.400 ;
        RECT 100.540 175.340 126.150 175.700 ;
        RECT 127.890 175.300 129.090 175.700 ;
        RECT 81.645 174.490 91.645 174.720 ;
        RECT 108.455 174.490 118.455 174.720 ;
        RECT 128.790 174.600 129.090 175.300 ;
        RECT 129.490 175.700 129.690 176.600 ;
        RECT 130.710 176.550 130.940 176.600 ;
        RECT 131.150 177.500 131.380 177.550 ;
        RECT 131.150 176.600 131.790 177.500 ;
        RECT 131.150 176.550 131.380 176.600 ;
        RECT 130.890 175.700 131.190 176.400 ;
        RECT 129.490 175.300 131.190 175.700 ;
        RECT 81.210 174.380 81.440 174.440 ;
        RECT 91.850 174.380 92.080 174.440 ;
        RECT 108.020 174.380 108.250 174.440 ;
        RECT 118.660 174.380 118.890 174.440 ;
        RECT 128.610 174.400 128.840 174.405 ;
        RECT 81.140 173.540 81.500 174.380 ;
        RECT 91.780 173.540 92.140 174.380 ;
        RECT 107.950 173.540 108.310 174.380 ;
        RECT 118.590 173.540 118.950 174.380 ;
        RECT 81.210 173.480 81.440 173.540 ;
        RECT 91.850 173.480 92.080 173.540 ;
        RECT 108.020 173.480 108.250 173.540 ;
        RECT 118.660 173.480 118.890 173.540 ;
        RECT 81.655 173.430 91.635 173.460 ;
        RECT 108.465 173.430 118.445 173.460 ;
        RECT 81.645 173.200 91.645 173.430 ;
        RECT 108.455 173.200 118.455 173.430 ;
        RECT 128.090 172.500 128.840 174.400 ;
        RECT 73.730 172.100 98.030 172.360 ;
        RECT 100.540 172.100 124.840 172.360 ;
        RECT 85.140 171.450 85.860 171.490 ;
        RECT 87.220 171.450 87.920 171.460 ;
        RECT 75.855 171.220 85.860 171.450 ;
        RECT 87.215 171.220 97.210 171.450 ;
        RECT 85.140 171.170 85.860 171.220 ;
        RECT 87.220 171.190 88.310 171.220 ;
        RECT 75.400 171.110 75.680 171.170 ;
        RECT 75.050 170.920 75.680 171.110 ;
        RECT 75.050 168.710 75.240 170.920 ;
        RECT 75.400 170.860 75.680 170.920 ;
        RECT 86.040 170.860 86.310 171.170 ;
        RECT 86.760 170.860 87.040 171.170 ;
        RECT 97.400 171.110 97.670 171.170 ;
        RECT 97.840 171.110 98.030 172.100 ;
        RECT 111.950 171.450 112.670 171.490 ;
        RECT 114.030 171.450 114.730 171.460 ;
        RECT 102.665 171.220 112.670 171.450 ;
        RECT 114.025 171.220 124.020 171.450 ;
        RECT 111.950 171.170 112.670 171.220 ;
        RECT 114.030 171.190 115.120 171.220 ;
        RECT 102.210 171.110 102.490 171.170 ;
        RECT 97.400 170.920 98.030 171.110 ;
        RECT 97.400 170.860 97.670 170.920 ;
        RECT 75.880 170.810 76.600 170.850 ;
        RECT 87.210 170.810 88.310 170.820 ;
        RECT 96.470 170.810 97.190 170.860 ;
        RECT 75.855 170.580 85.850 170.810 ;
        RECT 87.210 170.580 97.210 170.810 ;
        RECT 75.880 170.530 76.600 170.580 ;
        RECT 87.210 170.560 88.310 170.580 ;
        RECT 96.470 170.520 97.190 170.580 ;
        RECT 85.140 170.250 85.860 170.290 ;
        RECT 87.220 170.250 87.940 170.300 ;
        RECT 75.855 170.020 85.860 170.250 ;
        RECT 87.215 170.020 97.210 170.250 ;
        RECT 85.140 169.970 85.860 170.020 ;
        RECT 75.380 169.660 75.700 169.970 ;
        RECT 86.000 169.640 86.340 169.990 ;
        RECT 86.730 169.640 87.070 169.990 ;
        RECT 87.220 169.970 87.940 170.020 ;
        RECT 97.370 169.640 97.700 170.000 ;
        RECT 77.080 169.610 77.800 169.640 ;
        RECT 95.270 169.610 95.990 169.620 ;
        RECT 75.855 169.380 85.850 169.610 ;
        RECT 87.215 169.380 97.210 169.610 ;
        RECT 77.080 169.330 77.800 169.380 ;
        RECT 95.270 169.360 95.990 169.380 ;
        RECT 85.140 169.050 85.860 169.090 ;
        RECT 87.220 169.050 87.940 169.100 ;
        RECT 75.855 168.820 85.860 169.050 ;
        RECT 87.215 168.820 97.210 169.050 ;
        RECT 85.140 168.770 85.860 168.820 ;
        RECT 87.220 168.790 88.270 168.820 ;
        RECT 75.400 168.710 75.680 168.770 ;
        RECT 75.050 168.520 75.680 168.710 ;
        RECT 61.390 146.740 63.550 159.710 ;
        RECT 69.120 147.120 71.280 166.570 ;
        RECT 75.050 166.410 75.240 168.520 ;
        RECT 75.400 168.460 75.680 168.520 ;
        RECT 86.040 168.460 86.310 168.770 ;
        RECT 86.760 168.460 87.040 168.770 ;
        RECT 97.400 168.710 97.670 168.770 ;
        RECT 97.840 168.710 98.030 170.920 ;
        RECT 97.400 168.520 98.030 168.710 ;
        RECT 101.860 170.920 102.490 171.110 ;
        RECT 101.860 168.710 102.050 170.920 ;
        RECT 102.210 170.860 102.490 170.920 ;
        RECT 112.850 170.860 113.120 171.170 ;
        RECT 113.570 170.860 113.850 171.170 ;
        RECT 124.210 171.110 124.480 171.170 ;
        RECT 124.650 171.110 124.840 172.100 ;
        RECT 128.090 171.710 128.390 172.500 ;
        RECT 128.610 172.405 128.840 172.500 ;
        RECT 129.050 174.400 129.280 174.405 ;
        RECT 129.490 174.400 129.690 175.300 ;
        RECT 130.890 174.600 131.190 175.300 ;
        RECT 131.590 175.700 131.790 176.600 ;
        RECT 131.590 175.300 131.990 175.700 ;
        RECT 130.710 174.400 130.940 174.405 ;
        RECT 129.050 172.500 129.690 174.400 ;
        RECT 130.190 172.500 130.940 174.400 ;
        RECT 129.050 172.405 129.280 172.500 ;
        RECT 128.790 171.900 129.090 172.200 ;
        RECT 130.190 171.710 130.490 172.500 ;
        RECT 130.710 172.405 130.940 172.500 ;
        RECT 131.150 174.400 131.380 174.405 ;
        RECT 131.590 174.400 131.790 175.300 ;
        RECT 131.150 172.500 131.790 174.400 ;
        RECT 131.150 172.405 131.380 172.500 ;
        RECT 130.890 171.900 131.190 172.200 ;
        RECT 124.210 170.920 124.840 171.110 ;
        RECT 124.210 170.860 124.480 170.920 ;
        RECT 102.690 170.810 103.410 170.850 ;
        RECT 114.020 170.810 115.120 170.820 ;
        RECT 123.280 170.810 124.000 170.860 ;
        RECT 102.665 170.580 112.660 170.810 ;
        RECT 114.020 170.580 124.020 170.810 ;
        RECT 102.690 170.530 103.410 170.580 ;
        RECT 114.020 170.560 115.120 170.580 ;
        RECT 123.280 170.520 124.000 170.580 ;
        RECT 111.950 170.250 112.670 170.290 ;
        RECT 114.030 170.250 114.750 170.300 ;
        RECT 102.665 170.020 112.670 170.250 ;
        RECT 114.025 170.020 124.020 170.250 ;
        RECT 111.950 169.970 112.670 170.020 ;
        RECT 102.190 169.660 102.510 169.970 ;
        RECT 112.810 169.640 113.150 169.990 ;
        RECT 113.540 169.640 113.880 169.990 ;
        RECT 114.030 169.970 114.750 170.020 ;
        RECT 124.180 169.640 124.510 170.000 ;
        RECT 103.890 169.610 104.610 169.640 ;
        RECT 122.080 169.610 122.800 169.620 ;
        RECT 102.665 169.380 112.660 169.610 ;
        RECT 114.025 169.380 124.020 169.610 ;
        RECT 103.890 169.330 104.610 169.380 ;
        RECT 122.080 169.360 122.800 169.380 ;
        RECT 111.950 169.050 112.670 169.090 ;
        RECT 114.030 169.050 114.750 169.100 ;
        RECT 102.665 168.820 112.670 169.050 ;
        RECT 114.025 168.820 124.020 169.050 ;
        RECT 111.950 168.770 112.670 168.820 ;
        RECT 114.030 168.790 115.080 168.820 ;
        RECT 102.210 168.710 102.490 168.770 ;
        RECT 101.860 168.520 102.490 168.710 ;
        RECT 97.400 168.460 97.670 168.520 ;
        RECT 75.880 168.410 76.600 168.450 ;
        RECT 87.210 168.410 88.270 168.420 ;
        RECT 96.470 168.410 97.190 168.460 ;
        RECT 75.855 168.180 85.850 168.410 ;
        RECT 87.210 168.180 97.210 168.410 ;
        RECT 75.880 168.130 76.600 168.180 ;
        RECT 87.210 168.160 88.270 168.180 ;
        RECT 96.470 168.120 97.190 168.180 ;
        RECT 85.140 167.850 85.860 167.890 ;
        RECT 87.220 167.850 87.940 167.900 ;
        RECT 75.855 167.620 85.860 167.850 ;
        RECT 87.215 167.620 97.210 167.850 ;
        RECT 85.140 167.570 85.860 167.620 ;
        RECT 75.380 167.260 75.700 167.570 ;
        RECT 86.000 167.240 86.340 167.590 ;
        RECT 86.730 167.240 87.070 167.590 ;
        RECT 87.220 167.570 87.940 167.620 ;
        RECT 97.370 167.240 97.700 167.600 ;
        RECT 77.080 167.210 77.800 167.240 ;
        RECT 95.270 167.210 95.990 167.220 ;
        RECT 75.855 166.980 85.850 167.210 ;
        RECT 87.215 166.980 97.210 167.210 ;
        RECT 77.080 166.930 77.800 166.980 ;
        RECT 95.270 166.960 95.990 166.980 ;
        RECT 101.860 166.410 102.050 168.520 ;
        RECT 102.210 168.460 102.490 168.520 ;
        RECT 112.850 168.460 113.120 168.770 ;
        RECT 113.570 168.460 113.850 168.770 ;
        RECT 124.210 168.710 124.480 168.770 ;
        RECT 124.650 168.710 124.840 170.920 ;
        RECT 127.890 170.910 146.850 171.710 ;
        RECT 124.210 168.520 124.840 168.710 ;
        RECT 128.090 170.120 128.390 170.910 ;
        RECT 128.790 170.420 129.090 170.720 ;
        RECT 128.610 170.120 128.840 170.215 ;
        RECT 124.210 168.460 124.480 168.520 ;
        RECT 102.690 168.410 103.410 168.450 ;
        RECT 114.020 168.410 115.080 168.420 ;
        RECT 123.280 168.410 124.000 168.460 ;
        RECT 102.665 168.180 112.660 168.410 ;
        RECT 114.020 168.180 124.020 168.410 ;
        RECT 128.090 168.220 128.840 170.120 ;
        RECT 128.610 168.215 128.840 168.220 ;
        RECT 129.050 170.120 129.280 170.215 ;
        RECT 130.190 170.120 130.490 170.910 ;
        RECT 130.890 170.420 131.190 170.720 ;
        RECT 130.710 170.120 130.940 170.215 ;
        RECT 129.050 168.220 129.690 170.120 ;
        RECT 130.190 168.220 130.940 170.120 ;
        RECT 129.050 168.215 129.280 168.220 ;
        RECT 102.690 168.130 103.410 168.180 ;
        RECT 114.020 168.160 115.080 168.180 ;
        RECT 123.280 168.120 124.000 168.180 ;
        RECT 111.950 167.850 112.670 167.890 ;
        RECT 114.030 167.850 114.750 167.900 ;
        RECT 102.665 167.620 112.670 167.850 ;
        RECT 114.025 167.620 124.020 167.850 ;
        RECT 111.950 167.570 112.670 167.620 ;
        RECT 102.190 167.260 102.510 167.570 ;
        RECT 112.810 167.240 113.150 167.590 ;
        RECT 113.540 167.240 113.880 167.590 ;
        RECT 114.030 167.570 114.750 167.620 ;
        RECT 124.180 167.240 124.510 167.600 ;
        RECT 128.790 167.320 129.090 168.020 ;
        RECT 103.890 167.210 104.610 167.240 ;
        RECT 122.080 167.210 122.800 167.220 ;
        RECT 102.665 166.980 112.660 167.210 ;
        RECT 114.025 166.980 124.020 167.210 ;
        RECT 103.890 166.930 104.610 166.980 ;
        RECT 122.080 166.960 122.800 166.980 ;
        RECT 127.890 166.920 129.090 167.320 ;
        RECT 73.730 166.150 97.700 166.410 ;
        RECT 100.540 166.150 124.510 166.410 ;
        RECT 128.790 166.220 129.090 166.920 ;
        RECT 129.490 167.320 129.690 168.220 ;
        RECT 130.710 168.215 130.940 168.220 ;
        RECT 131.150 170.120 131.380 170.215 ;
        RECT 131.150 168.220 131.790 170.120 ;
        RECT 131.150 168.215 131.380 168.220 ;
        RECT 130.890 167.320 131.190 168.020 ;
        RECT 129.490 166.920 131.190 167.320 ;
        RECT 128.610 166.020 128.840 166.070 ;
        RECT 77.070 165.750 97.190 166.010 ;
        RECT 103.880 165.750 124.000 166.010 ;
        RECT 75.870 165.350 95.990 165.610 ;
        RECT 102.680 165.350 122.800 165.610 ;
        RECT 128.090 165.120 128.840 166.020 ;
        RECT 74.390 164.470 78.770 164.490 ;
        RECT 80.640 164.470 85.620 164.490 ;
        RECT 87.610 164.470 92.590 164.490 ;
        RECT 74.390 164.230 79.170 164.470 ;
        RECT 80.630 164.240 85.630 164.470 ;
        RECT 87.600 164.240 92.600 164.470 ;
        RECT 80.640 164.230 85.620 164.240 ;
        RECT 87.610 164.230 92.590 164.240 ;
        RECT 93.930 164.230 98.680 164.490 ;
        RECT 74.390 163.840 74.620 164.230 ;
        RECT 78.940 164.130 79.170 164.230 ;
        RECT 93.930 164.210 94.290 164.230 ;
        RECT 93.930 164.190 94.130 164.210 ;
        RECT 80.240 164.130 80.470 164.190 ;
        RECT 85.790 164.130 86.020 164.190 ;
        RECT 87.210 164.130 87.440 164.190 ;
        RECT 92.760 164.130 92.990 164.190 ;
        RECT 93.900 164.130 94.130 164.190 ;
        RECT 78.940 163.840 80.470 164.130 ;
        RECT 85.720 163.840 86.080 164.130 ;
        RECT 74.390 163.580 86.080 163.840 ;
        RECT 74.390 163.230 74.620 163.580 ;
        RECT 78.940 163.290 80.470 163.580 ;
        RECT 85.720 163.290 86.080 163.580 ;
        RECT 87.150 163.840 87.510 164.130 ;
        RECT 92.760 163.840 94.130 164.130 ;
        RECT 98.450 163.840 98.680 164.230 ;
        RECT 87.150 163.580 98.680 163.840 ;
        RECT 87.150 163.290 87.510 163.580 ;
        RECT 92.760 163.290 94.130 163.580 ;
        RECT 78.940 163.230 79.170 163.290 ;
        RECT 80.240 163.230 80.470 163.290 ;
        RECT 85.790 163.230 86.020 163.290 ;
        RECT 87.210 163.230 87.440 163.290 ;
        RECT 92.760 163.230 92.990 163.290 ;
        RECT 93.900 163.230 94.130 163.290 ;
        RECT 98.450 163.230 98.680 163.580 ;
        RECT 101.200 164.470 105.580 164.490 ;
        RECT 107.450 164.470 112.430 164.490 ;
        RECT 114.420 164.470 119.400 164.490 ;
        RECT 101.200 164.230 105.980 164.470 ;
        RECT 107.440 164.240 112.440 164.470 ;
        RECT 114.410 164.240 119.410 164.470 ;
        RECT 107.450 164.230 112.430 164.240 ;
        RECT 114.420 164.230 119.400 164.240 ;
        RECT 120.740 164.230 125.490 164.490 ;
        RECT 128.090 164.420 128.390 165.120 ;
        RECT 128.610 165.070 128.840 165.120 ;
        RECT 129.050 166.020 129.280 166.070 ;
        RECT 129.490 166.020 129.690 166.920 ;
        RECT 130.890 166.220 131.190 166.920 ;
        RECT 131.590 167.320 131.790 168.220 ;
        RECT 131.590 166.920 131.990 167.320 ;
        RECT 130.710 166.020 130.940 166.070 ;
        RECT 129.050 165.120 129.690 166.020 ;
        RECT 130.190 165.120 130.940 166.020 ;
        RECT 129.050 165.070 129.280 165.120 ;
        RECT 128.790 164.620 129.090 164.920 ;
        RECT 130.190 164.420 130.490 165.120 ;
        RECT 130.710 165.070 130.940 165.120 ;
        RECT 131.150 166.020 131.380 166.070 ;
        RECT 131.590 166.020 131.790 166.920 ;
        RECT 131.150 165.120 131.790 166.020 ;
        RECT 131.150 165.070 131.380 165.120 ;
        RECT 130.890 164.620 131.190 164.920 ;
        RECT 101.200 163.840 101.430 164.230 ;
        RECT 105.750 164.130 105.980 164.230 ;
        RECT 120.740 164.210 121.100 164.230 ;
        RECT 120.740 164.190 120.940 164.210 ;
        RECT 107.050 164.130 107.280 164.190 ;
        RECT 112.600 164.130 112.830 164.190 ;
        RECT 114.020 164.130 114.250 164.190 ;
        RECT 119.570 164.130 119.800 164.190 ;
        RECT 120.710 164.130 120.940 164.190 ;
        RECT 105.750 163.840 107.280 164.130 ;
        RECT 112.530 163.840 112.890 164.130 ;
        RECT 101.200 163.580 112.890 163.840 ;
        RECT 101.200 163.230 101.430 163.580 ;
        RECT 105.750 163.290 107.280 163.580 ;
        RECT 112.530 163.290 112.890 163.580 ;
        RECT 113.960 163.840 114.320 164.130 ;
        RECT 119.570 163.840 120.940 164.130 ;
        RECT 125.260 163.840 125.490 164.230 ;
        RECT 127.890 164.020 146.850 164.420 ;
        RECT 113.960 163.580 125.490 163.840 ;
        RECT 113.960 163.290 114.320 163.580 ;
        RECT 119.570 163.290 120.940 163.580 ;
        RECT 105.750 163.230 105.980 163.290 ;
        RECT 107.050 163.230 107.280 163.290 ;
        RECT 112.600 163.230 112.830 163.290 ;
        RECT 114.020 163.230 114.250 163.290 ;
        RECT 119.570 163.230 119.800 163.290 ;
        RECT 120.710 163.230 120.940 163.290 ;
        RECT 125.260 163.230 125.490 163.580 ;
        RECT 74.780 162.950 78.780 163.180 ;
        RECT 80.630 162.950 85.630 163.180 ;
        RECT 87.600 162.950 92.600 163.180 ;
        RECT 94.290 162.950 98.290 163.180 ;
        RECT 101.590 162.950 105.590 163.180 ;
        RECT 107.440 162.950 112.440 163.180 ;
        RECT 114.410 162.950 119.410 163.180 ;
        RECT 121.100 162.950 125.100 163.180 ;
        RECT 75.090 162.580 78.460 162.950 ;
        RECT 81.380 162.580 84.750 162.950 ;
        RECT 88.490 162.580 91.860 162.950 ;
        RECT 101.900 162.580 105.270 162.950 ;
        RECT 108.190 162.580 111.560 162.950 ;
        RECT 115.300 162.580 118.670 162.950 ;
        RECT 73.730 162.410 99.340 162.580 ;
        RECT 73.730 160.180 79.650 162.410 ;
        RECT 80.640 162.040 85.620 162.060 ;
        RECT 87.610 162.040 92.590 162.060 ;
        RECT 80.630 161.810 85.630 162.040 ;
        RECT 87.600 161.810 92.600 162.040 ;
        RECT 80.640 161.800 85.620 161.810 ;
        RECT 87.610 161.800 92.590 161.810 ;
        RECT 80.240 161.420 80.470 161.760 ;
        RECT 85.790 161.700 86.020 161.760 ;
        RECT 87.210 161.700 87.440 161.760 ;
        RECT 85.720 161.420 86.080 161.700 ;
        RECT 80.240 161.160 86.080 161.420 ;
        RECT 80.240 160.800 80.470 161.160 ;
        RECT 85.720 160.860 86.080 161.160 ;
        RECT 87.150 161.420 87.510 161.700 ;
        RECT 92.760 161.420 92.990 161.760 ;
        RECT 87.150 161.160 92.990 161.420 ;
        RECT 87.150 160.860 87.510 161.160 ;
        RECT 85.790 160.800 86.020 160.860 ;
        RECT 87.210 160.800 87.440 160.860 ;
        RECT 92.760 160.800 92.990 161.160 ;
        RECT 80.630 160.520 85.630 160.750 ;
        RECT 87.600 160.520 92.600 160.750 ;
        RECT 80.690 160.180 85.570 160.520 ;
        RECT 87.660 160.180 92.540 160.520 ;
        RECT 93.420 160.180 99.340 162.410 ;
        RECT 73.730 159.800 99.340 160.180 ;
        RECT 100.540 162.410 126.150 162.580 ;
        RECT 100.540 160.180 106.460 162.410 ;
        RECT 107.450 162.040 112.430 162.060 ;
        RECT 114.420 162.040 119.400 162.060 ;
        RECT 107.440 161.810 112.440 162.040 ;
        RECT 114.410 161.810 119.410 162.040 ;
        RECT 107.450 161.800 112.430 161.810 ;
        RECT 114.420 161.800 119.400 161.810 ;
        RECT 107.050 161.420 107.280 161.760 ;
        RECT 112.600 161.700 112.830 161.760 ;
        RECT 114.020 161.700 114.250 161.760 ;
        RECT 112.530 161.420 112.890 161.700 ;
        RECT 107.050 161.160 112.890 161.420 ;
        RECT 107.050 160.800 107.280 161.160 ;
        RECT 112.530 160.860 112.890 161.160 ;
        RECT 113.960 161.420 114.320 161.700 ;
        RECT 119.570 161.420 119.800 161.760 ;
        RECT 113.960 161.160 119.800 161.420 ;
        RECT 113.960 160.860 114.320 161.160 ;
        RECT 112.600 160.800 112.830 160.860 ;
        RECT 114.020 160.800 114.250 160.860 ;
        RECT 119.570 160.800 119.800 161.160 ;
        RECT 107.440 160.520 112.440 160.750 ;
        RECT 114.410 160.520 119.410 160.750 ;
        RECT 107.500 160.180 112.380 160.520 ;
        RECT 114.470 160.180 119.350 160.520 ;
        RECT 120.230 160.180 126.150 162.410 ;
        RECT 100.540 159.800 126.150 160.180 ;
        RECT 93.420 159.790 99.340 159.800 ;
        RECT 100.530 159.790 126.150 159.800 ;
        RECT 100.530 159.420 126.140 159.790 ;
        RECT 100.530 157.190 106.450 159.420 ;
        RECT 107.490 159.080 112.370 159.420 ;
        RECT 114.460 159.080 119.340 159.420 ;
        RECT 107.430 158.850 112.430 159.080 ;
        RECT 114.400 158.850 119.400 159.080 ;
        RECT 107.040 158.440 107.270 158.800 ;
        RECT 112.590 158.740 112.820 158.800 ;
        RECT 114.010 158.740 114.240 158.800 ;
        RECT 112.520 158.440 112.880 158.740 ;
        RECT 107.040 158.180 112.880 158.440 ;
        RECT 107.040 157.840 107.270 158.180 ;
        RECT 112.520 157.900 112.880 158.180 ;
        RECT 113.950 158.440 114.310 158.740 ;
        RECT 119.560 158.440 119.790 158.800 ;
        RECT 113.950 158.180 119.790 158.440 ;
        RECT 113.950 157.900 114.310 158.180 ;
        RECT 112.590 157.840 112.820 157.900 ;
        RECT 114.010 157.840 114.240 157.900 ;
        RECT 119.560 157.840 119.790 158.180 ;
        RECT 107.440 157.790 112.420 157.800 ;
        RECT 114.410 157.790 119.390 157.800 ;
        RECT 107.430 157.560 112.430 157.790 ;
        RECT 114.400 157.560 119.400 157.790 ;
        RECT 107.440 157.540 112.420 157.560 ;
        RECT 114.410 157.540 119.390 157.560 ;
        RECT 120.220 157.190 126.140 159.420 ;
        RECT 100.530 157.020 126.140 157.190 ;
        RECT 101.890 156.650 105.260 157.020 ;
        RECT 108.180 156.650 111.550 157.020 ;
        RECT 115.290 156.650 118.660 157.020 ;
        RECT 101.580 156.420 105.580 156.650 ;
        RECT 107.430 156.420 112.430 156.650 ;
        RECT 114.400 156.420 119.400 156.650 ;
        RECT 121.090 156.420 125.090 156.650 ;
        RECT 101.190 156.020 101.420 156.370 ;
        RECT 105.740 156.310 105.970 156.370 ;
        RECT 107.040 156.310 107.270 156.370 ;
        RECT 112.590 156.310 112.820 156.370 ;
        RECT 114.010 156.310 114.240 156.370 ;
        RECT 119.560 156.310 119.790 156.370 ;
        RECT 120.700 156.310 120.930 156.370 ;
        RECT 105.740 156.020 107.270 156.310 ;
        RECT 112.520 156.020 112.880 156.310 ;
        RECT 101.190 155.760 112.880 156.020 ;
        RECT 101.190 155.370 101.420 155.760 ;
        RECT 105.740 155.470 107.270 155.760 ;
        RECT 112.520 155.470 112.880 155.760 ;
        RECT 113.950 156.020 114.310 156.310 ;
        RECT 119.560 156.020 120.930 156.310 ;
        RECT 125.250 156.020 125.480 156.370 ;
        RECT 113.950 155.760 125.480 156.020 ;
        RECT 113.950 155.470 114.310 155.760 ;
        RECT 119.560 155.470 120.930 155.760 ;
        RECT 105.740 155.370 105.970 155.470 ;
        RECT 107.040 155.410 107.270 155.470 ;
        RECT 112.590 155.410 112.820 155.470 ;
        RECT 114.010 155.410 114.240 155.470 ;
        RECT 119.560 155.410 119.790 155.470 ;
        RECT 120.700 155.410 120.930 155.470 ;
        RECT 120.730 155.390 120.930 155.410 ;
        RECT 120.730 155.370 121.090 155.390 ;
        RECT 125.250 155.370 125.480 155.760 ;
        RECT 101.190 155.130 105.970 155.370 ;
        RECT 107.440 155.360 112.420 155.370 ;
        RECT 114.410 155.360 119.390 155.370 ;
        RECT 107.430 155.130 112.430 155.360 ;
        RECT 114.400 155.130 119.400 155.360 ;
        RECT 101.190 155.110 105.570 155.130 ;
        RECT 107.440 155.110 112.420 155.130 ;
        RECT 114.410 155.110 119.390 155.130 ;
        RECT 120.730 155.110 125.480 155.370 ;
        RECT 84.010 153.300 84.390 154.400 ;
        RECT 85.070 153.750 89.120 153.800 ;
        RECT 85.010 153.520 89.120 153.750 ;
        RECT 85.070 153.500 89.120 153.520 ;
        RECT 86.040 153.360 89.120 153.500 ;
        RECT 84.730 153.300 84.960 153.360 ;
        RECT 84.010 148.420 84.960 153.300 ;
        RECT 84.010 147.310 84.390 148.420 ;
        RECT 84.730 148.360 84.960 148.420 ;
        RECT 86.020 151.420 89.120 153.360 ;
        RECT 90.250 151.420 94.200 153.580 ;
        RECT 95.330 153.490 99.470 153.580 ;
        RECT 95.330 153.260 99.530 153.490 ;
        RECT 100.150 153.450 100.530 154.410 ;
        RECT 102.670 153.990 122.790 154.250 ;
        RECT 103.870 153.590 123.990 153.850 ;
        RECT 95.330 153.230 99.470 153.260 ;
        RECT 95.330 153.055 98.490 153.230 ;
        RECT 100.150 153.190 124.500 153.450 ;
        RECT 95.330 151.420 98.520 153.055 ;
        RECT 86.020 148.360 86.250 151.420 ;
        RECT 85.010 147.970 85.990 148.200 ;
        RECT 85.070 147.310 85.990 147.970 ;
        RECT 60.560 146.290 72.110 146.740 ;
        RECT 87.710 142.420 91.660 144.580 ;
        RECT 92.790 142.420 96.740 144.580 ;
        RECT 98.290 143.055 98.520 151.420 ;
        RECT 99.580 153.010 99.810 153.055 ;
        RECT 100.150 153.010 100.530 153.190 ;
        RECT 99.580 147.500 100.530 153.010 ;
        RECT 101.850 151.080 102.040 153.190 ;
        RECT 103.880 152.620 104.600 152.670 ;
        RECT 122.070 152.620 122.790 152.640 ;
        RECT 102.655 152.390 112.650 152.620 ;
        RECT 114.015 152.390 124.010 152.620 ;
        RECT 103.880 152.360 104.600 152.390 ;
        RECT 122.070 152.380 122.790 152.390 ;
        RECT 102.180 152.030 102.500 152.340 ;
        RECT 111.940 151.980 112.660 152.030 ;
        RECT 112.800 152.010 113.140 152.360 ;
        RECT 113.530 152.010 113.870 152.360 ;
        RECT 114.020 151.980 114.740 152.030 ;
        RECT 124.170 152.000 124.500 152.360 ;
        RECT 102.655 151.750 112.660 151.980 ;
        RECT 114.015 151.750 124.010 151.980 ;
        RECT 111.940 151.710 112.660 151.750 ;
        RECT 114.020 151.700 114.740 151.750 ;
        RECT 102.680 151.420 103.400 151.470 ;
        RECT 114.010 151.420 115.070 151.440 ;
        RECT 123.270 151.420 123.990 151.480 ;
        RECT 102.655 151.190 112.650 151.420 ;
        RECT 114.010 151.190 124.010 151.420 ;
        RECT 102.680 151.150 103.400 151.190 ;
        RECT 114.010 151.180 115.070 151.190 ;
        RECT 123.270 151.140 123.990 151.190 ;
        RECT 102.200 151.080 102.480 151.140 ;
        RECT 101.850 150.890 102.480 151.080 ;
        RECT 101.850 148.680 102.040 150.890 ;
        RECT 102.200 150.830 102.480 150.890 ;
        RECT 112.840 150.830 113.110 151.140 ;
        RECT 113.560 150.830 113.840 151.140 ;
        RECT 124.200 151.080 124.470 151.140 ;
        RECT 124.200 150.890 124.830 151.080 ;
        RECT 124.200 150.830 124.470 150.890 ;
        RECT 111.940 150.780 112.660 150.830 ;
        RECT 114.020 150.780 115.070 150.810 ;
        RECT 102.655 150.550 112.660 150.780 ;
        RECT 114.015 150.550 124.010 150.780 ;
        RECT 111.940 150.510 112.660 150.550 ;
        RECT 114.020 150.500 114.740 150.550 ;
        RECT 103.880 150.220 104.600 150.270 ;
        RECT 122.070 150.220 122.790 150.240 ;
        RECT 102.655 149.990 112.650 150.220 ;
        RECT 114.015 149.990 124.010 150.220 ;
        RECT 103.880 149.960 104.600 149.990 ;
        RECT 122.070 149.980 122.790 149.990 ;
        RECT 102.180 149.630 102.500 149.940 ;
        RECT 111.940 149.580 112.660 149.630 ;
        RECT 112.800 149.610 113.140 149.960 ;
        RECT 113.530 149.610 113.870 149.960 ;
        RECT 114.020 149.580 114.740 149.630 ;
        RECT 124.170 149.600 124.500 149.960 ;
        RECT 102.655 149.350 112.660 149.580 ;
        RECT 114.015 149.350 124.010 149.580 ;
        RECT 111.940 149.310 112.660 149.350 ;
        RECT 114.020 149.300 114.740 149.350 ;
        RECT 102.680 149.020 103.400 149.070 ;
        RECT 114.010 149.020 115.110 149.040 ;
        RECT 123.270 149.020 123.990 149.080 ;
        RECT 102.655 148.790 112.650 149.020 ;
        RECT 114.010 148.790 124.010 149.020 ;
        RECT 102.680 148.750 103.400 148.790 ;
        RECT 114.010 148.780 115.110 148.790 ;
        RECT 123.270 148.740 123.990 148.790 ;
        RECT 102.200 148.680 102.480 148.740 ;
        RECT 101.850 148.490 102.480 148.680 ;
        RECT 102.200 148.430 102.480 148.490 ;
        RECT 112.840 148.430 113.110 148.740 ;
        RECT 113.560 148.430 113.840 148.740 ;
        RECT 124.200 148.680 124.470 148.740 ;
        RECT 124.640 148.680 124.830 150.890 ;
        RECT 124.200 148.490 124.830 148.680 ;
        RECT 124.200 148.430 124.470 148.490 ;
        RECT 111.940 148.380 112.660 148.430 ;
        RECT 114.020 148.380 115.110 148.410 ;
        RECT 102.655 148.150 112.660 148.380 ;
        RECT 114.015 148.150 124.010 148.380 ;
        RECT 111.940 148.110 112.660 148.150 ;
        RECT 114.020 148.140 114.720 148.150 ;
        RECT 124.640 147.500 124.830 148.490 ;
        RECT 99.580 147.240 124.830 147.500 ;
        RECT 99.580 144.260 100.530 147.240 ;
        RECT 108.445 146.170 118.445 146.400 ;
        RECT 108.455 146.140 118.435 146.170 ;
        RECT 108.010 146.060 108.240 146.120 ;
        RECT 118.650 146.060 118.880 146.120 ;
        RECT 107.940 145.220 108.300 146.060 ;
        RECT 118.580 145.220 118.940 146.060 ;
        RECT 108.010 145.160 108.240 145.220 ;
        RECT 118.650 145.160 118.880 145.220 ;
        RECT 108.445 144.880 118.445 145.110 ;
        RECT 99.580 143.900 126.140 144.260 ;
        RECT 99.580 143.100 103.770 143.900 ;
        RECT 99.580 143.055 99.810 143.100 ;
        RECT 98.550 142.850 99.470 142.910 ;
        RECT 98.550 142.620 99.530 142.850 ;
        RECT 98.550 142.140 99.470 142.620 ;
        RECT 100.150 141.670 103.770 143.100 ;
        RECT 104.070 143.280 112.940 143.540 ;
        RECT 114.170 143.530 122.150 143.540 ;
        RECT 114.165 143.300 122.165 143.530 ;
        RECT 114.170 143.280 122.150 143.300 ;
        RECT 104.070 142.890 104.300 143.280 ;
        RECT 112.710 143.190 112.940 143.280 ;
        RECT 113.730 143.190 113.960 143.250 ;
        RECT 112.710 142.890 113.960 143.190 ;
        RECT 122.370 142.890 122.600 143.250 ;
        RECT 104.070 142.630 122.600 142.890 ;
        RECT 104.070 142.290 104.300 142.630 ;
        RECT 112.710 142.350 113.960 142.630 ;
        RECT 112.710 142.290 112.940 142.350 ;
        RECT 113.730 142.290 113.960 142.350 ;
        RECT 122.370 142.290 122.600 142.630 ;
        RECT 104.505 142.010 112.505 142.240 ;
        RECT 114.165 142.010 122.165 142.240 ;
        RECT 104.565 141.670 112.445 142.010 ;
        RECT 114.225 141.670 122.105 142.010 ;
        RECT 122.900 141.670 126.140 143.900 ;
        RECT 100.150 141.590 126.140 141.670 ;
        RECT 100.530 141.290 126.140 141.590 ;
      LAYER met2 ;
        RECT 73.730 214.640 86.660 214.900 ;
        RECT 100.540 214.640 113.470 214.900 ;
        RECT 127.890 214.650 146.850 215.050 ;
        RECT 77.760 213.340 85.640 213.390 ;
        RECT 73.860 213.080 85.640 213.340 ;
        RECT 73.860 199.080 74.120 213.080 ;
        RECT 77.760 213.030 85.640 213.080 ;
        RECT 81.190 211.110 81.450 211.450 ;
        RECT 86.400 211.110 86.660 214.640 ;
        RECT 87.420 213.340 95.300 213.390 ;
        RECT 104.570 213.340 112.450 213.390 ;
        RECT 87.420 213.080 99.340 213.340 ;
        RECT 100.670 213.080 112.450 213.340 ;
        RECT 87.420 213.030 95.300 213.080 ;
        RECT 91.830 211.110 92.090 211.450 ;
        RECT 81.190 210.850 92.090 211.110 ;
        RECT 81.190 210.510 81.450 210.850 ;
        RECT 86.400 210.840 86.660 210.850 ;
        RECT 81.705 210.170 91.585 210.530 ;
        RECT 91.830 210.510 92.090 210.850 ;
        RECT 85.130 209.685 87.940 210.170 ;
        RECT 75.370 206.660 75.710 209.380 ;
        RECT 75.370 204.610 75.700 206.660 ;
        RECT 75.370 204.260 75.710 204.610 ;
        RECT 75.880 201.560 76.600 207.870 ;
        RECT 77.080 202.700 77.800 206.660 ;
        RECT 85.140 204.610 85.860 209.685 ;
        RECT 86.000 204.260 86.340 209.380 ;
        RECT 86.730 203.170 87.070 207.010 ;
        RECT 87.220 204.590 87.940 209.685 ;
        RECT 77.540 201.980 77.800 202.700 ;
        RECT 95.270 202.370 95.990 206.640 ;
        RECT 95.270 202.320 95.940 202.370 ;
        RECT 80.690 201.980 80.950 201.990 ;
        RECT 95.270 201.980 95.530 202.320 ;
        RECT 77.540 201.720 80.950 201.980 ;
        RECT 80.690 201.560 80.950 201.720 ;
        RECT 92.280 201.720 95.530 201.980 ;
        RECT 92.280 201.560 92.540 201.720 ;
        RECT 96.470 201.560 97.190 207.880 ;
        RECT 97.370 203.170 97.700 207.020 ;
        RECT 74.840 201.200 78.720 201.560 ;
        RECT 80.690 201.200 85.570 201.560 ;
        RECT 87.660 201.200 92.540 201.560 ;
        RECT 94.340 201.200 98.220 201.560 ;
        RECT 80.690 199.080 85.570 199.130 ;
        RECT 73.860 198.820 85.570 199.080 ;
        RECT 80.690 198.770 85.570 198.820 ;
        RECT 85.770 197.830 86.030 201.200 ;
        RECT 87.200 197.830 87.460 201.200 ;
        RECT 87.660 199.080 92.540 199.130 ;
        RECT 98.950 199.080 99.210 213.080 ;
        RECT 87.660 198.820 99.210 199.080 ;
        RECT 100.670 199.080 100.930 213.080 ;
        RECT 104.570 213.030 112.450 213.080 ;
        RECT 108.000 211.110 108.260 211.450 ;
        RECT 113.210 211.110 113.470 214.640 ;
        RECT 114.230 213.340 122.110 213.390 ;
        RECT 114.230 213.080 126.150 213.340 ;
        RECT 114.230 213.030 122.110 213.080 ;
        RECT 118.640 211.110 118.900 211.450 ;
        RECT 108.000 210.850 118.900 211.110 ;
        RECT 108.000 210.510 108.260 210.850 ;
        RECT 113.210 210.840 113.470 210.850 ;
        RECT 108.515 210.170 118.395 210.530 ;
        RECT 118.640 210.510 118.900 210.850 ;
        RECT 111.940 209.685 114.750 210.170 ;
        RECT 102.180 206.660 102.520 209.380 ;
        RECT 102.180 204.610 102.510 206.660 ;
        RECT 102.180 204.260 102.520 204.610 ;
        RECT 102.690 201.560 103.410 207.870 ;
        RECT 103.890 202.700 104.610 206.660 ;
        RECT 111.950 204.610 112.670 209.685 ;
        RECT 112.810 204.260 113.150 209.380 ;
        RECT 113.540 203.170 113.880 207.010 ;
        RECT 114.030 204.590 114.750 209.685 ;
        RECT 104.350 201.980 104.610 202.700 ;
        RECT 122.080 202.370 122.800 206.640 ;
        RECT 122.080 202.320 122.750 202.370 ;
        RECT 107.500 201.980 107.760 201.990 ;
        RECT 122.080 201.980 122.340 202.320 ;
        RECT 104.350 201.720 107.760 201.980 ;
        RECT 107.500 201.560 107.760 201.720 ;
        RECT 119.090 201.720 122.340 201.980 ;
        RECT 119.090 201.560 119.350 201.720 ;
        RECT 123.280 201.560 124.000 207.880 ;
        RECT 124.180 203.170 124.510 207.020 ;
        RECT 101.650 201.200 105.530 201.560 ;
        RECT 107.500 201.200 112.380 201.560 ;
        RECT 114.470 201.200 119.350 201.560 ;
        RECT 121.150 201.200 125.030 201.560 ;
        RECT 107.500 199.080 112.380 199.130 ;
        RECT 100.670 198.820 112.380 199.080 ;
        RECT 87.660 198.770 92.540 198.820 ;
        RECT 107.500 198.770 112.380 198.820 ;
        RECT 112.580 197.830 112.840 201.200 ;
        RECT 114.010 197.830 114.270 201.200 ;
        RECT 114.470 199.080 119.350 199.130 ;
        RECT 125.760 199.080 126.020 213.080 ;
        RECT 131.240 212.840 131.670 213.800 ;
        RECT 134.140 212.840 134.540 213.840 ;
        RECT 131.240 212.480 134.540 212.840 ;
        RECT 136.560 212.490 136.950 213.750 ;
        RECT 131.240 212.050 131.670 212.480 ;
        RECT 134.140 212.110 134.540 212.480 ;
        RECT 135.240 211.810 139.770 212.210 ;
        RECT 135.240 211.550 135.810 211.810 ;
        RECT 132.990 209.980 133.320 210.920 ;
        RECT 133.610 210.700 136.500 211.030 ;
        RECT 140.580 210.690 143.760 211.070 ;
        RECT 132.940 208.330 136.520 208.620 ;
        RECT 127.890 207.360 146.850 208.160 ;
        RECT 132.940 206.900 136.520 207.190 ;
        RECT 138.210 206.900 141.790 207.190 ;
        RECT 139.370 205.860 139.770 206.560 ;
        RECT 133.000 205.450 133.310 205.470 ;
        RECT 132.950 203.780 133.350 205.450 ;
        RECT 133.610 204.490 136.500 204.820 ;
        RECT 138.260 204.020 138.590 205.540 ;
        RECT 140.580 205.300 141.020 206.550 ;
        RECT 141.840 205.840 142.230 206.590 ;
        RECT 138.880 204.490 141.770 204.820 ;
        RECT 142.840 204.460 143.840 204.860 ;
        RECT 142.840 204.020 143.120 204.460 ;
        RECT 135.290 203.690 143.120 204.020 ;
        RECT 131.250 202.830 131.680 203.460 ;
        RECT 134.120 202.830 134.550 203.440 ;
        RECT 135.290 203.210 135.760 203.690 ;
        RECT 131.250 202.430 134.550 202.830 ;
        RECT 131.250 201.720 131.680 202.430 ;
        RECT 134.120 201.700 134.550 202.430 ;
        RECT 136.530 201.880 136.980 203.310 ;
        RECT 127.890 200.070 146.850 200.870 ;
        RECT 114.470 198.820 126.020 199.080 ;
        RECT 114.470 198.770 119.350 198.820 ;
        RECT 135.220 198.680 142.220 199.180 ;
        RECT 131.270 197.830 131.710 198.180 ;
        RECT 134.130 197.830 134.520 198.320 ;
        RECT 135.220 198.160 135.800 198.680 ;
        RECT 131.270 197.480 134.520 197.830 ;
        RECT 136.530 197.490 136.960 198.240 ;
        RECT 80.690 194.820 85.570 194.870 ;
        RECT 73.860 194.560 85.570 194.820 ;
        RECT 73.860 180.560 74.120 194.560 ;
        RECT 80.690 194.510 85.570 194.560 ;
        RECT 85.770 192.440 86.030 195.810 ;
        RECT 87.200 192.440 87.460 195.810 ;
        RECT 87.660 194.820 92.540 194.870 ;
        RECT 107.500 194.820 112.380 194.870 ;
        RECT 87.660 194.560 99.210 194.820 ;
        RECT 87.660 194.510 92.540 194.560 ;
        RECT 74.840 192.080 78.720 192.440 ;
        RECT 80.690 192.080 85.570 192.440 ;
        RECT 87.660 192.080 92.540 192.440 ;
        RECT 94.340 192.080 98.220 192.440 ;
        RECT 75.370 189.030 75.710 189.380 ;
        RECT 75.370 186.980 75.700 189.030 ;
        RECT 75.370 184.260 75.710 186.980 ;
        RECT 75.880 185.770 76.600 192.080 ;
        RECT 80.690 191.920 80.950 192.080 ;
        RECT 77.540 191.660 80.950 191.920 ;
        RECT 92.280 191.920 92.540 192.080 ;
        RECT 92.280 191.660 95.530 191.920 ;
        RECT 77.540 190.940 77.800 191.660 ;
        RECT 80.690 191.650 80.950 191.660 ;
        RECT 77.080 186.980 77.800 190.940 ;
        RECT 95.270 191.320 95.530 191.660 ;
        RECT 95.270 191.270 95.940 191.320 ;
        RECT 85.140 183.955 85.860 189.030 ;
        RECT 86.000 184.260 86.340 189.380 ;
        RECT 86.730 186.630 87.070 190.470 ;
        RECT 87.220 183.955 87.940 189.050 ;
        RECT 95.270 187.000 95.990 191.270 ;
        RECT 96.470 185.760 97.190 192.080 ;
        RECT 97.370 186.620 97.700 190.470 ;
        RECT 85.130 183.470 87.940 183.955 ;
        RECT 81.190 182.790 81.450 183.130 ;
        RECT 81.705 183.110 91.585 183.470 ;
        RECT 86.400 182.790 86.660 182.800 ;
        RECT 91.830 182.790 92.090 183.130 ;
        RECT 81.190 182.530 92.090 182.790 ;
        RECT 81.190 182.190 81.450 182.530 ;
        RECT 77.760 180.560 85.640 180.610 ;
        RECT 73.860 180.300 85.640 180.560 ;
        RECT 77.760 180.250 85.640 180.300 ;
        RECT 86.400 179.000 86.660 182.530 ;
        RECT 91.830 182.190 92.090 182.530 ;
        RECT 87.420 180.560 95.300 180.610 ;
        RECT 98.950 180.560 99.210 194.560 ;
        RECT 100.670 194.560 112.380 194.820 ;
        RECT 100.670 180.560 100.930 194.560 ;
        RECT 107.500 194.510 112.380 194.560 ;
        RECT 112.580 192.440 112.840 195.810 ;
        RECT 114.010 192.440 114.270 195.810 ;
        RECT 132.990 195.060 133.320 197.160 ;
        RECT 133.610 196.120 136.500 196.450 ;
        RECT 141.430 195.620 142.110 196.570 ;
        RECT 141.430 195.060 141.760 195.620 ;
        RECT 114.470 194.820 119.350 194.870 ;
        RECT 114.470 194.560 126.020 194.820 ;
        RECT 132.990 194.720 141.760 195.060 ;
        RECT 114.470 194.510 119.350 194.560 ;
        RECT 101.650 192.080 105.530 192.440 ;
        RECT 107.500 192.080 112.380 192.440 ;
        RECT 114.470 192.080 119.350 192.440 ;
        RECT 121.150 192.080 125.030 192.440 ;
        RECT 102.180 189.030 102.520 189.380 ;
        RECT 102.180 186.980 102.510 189.030 ;
        RECT 102.180 184.260 102.520 186.980 ;
        RECT 102.690 185.770 103.410 192.080 ;
        RECT 107.500 191.920 107.760 192.080 ;
        RECT 104.350 191.660 107.760 191.920 ;
        RECT 119.090 191.920 119.350 192.080 ;
        RECT 119.090 191.660 122.340 191.920 ;
        RECT 104.350 190.940 104.610 191.660 ;
        RECT 107.500 191.650 107.760 191.660 ;
        RECT 103.890 186.980 104.610 190.940 ;
        RECT 122.080 191.320 122.340 191.660 ;
        RECT 122.080 191.270 122.750 191.320 ;
        RECT 111.950 183.955 112.670 189.030 ;
        RECT 112.810 184.260 113.150 189.380 ;
        RECT 113.540 186.630 113.880 190.470 ;
        RECT 114.030 183.955 114.750 189.050 ;
        RECT 122.080 187.000 122.800 191.270 ;
        RECT 123.280 185.760 124.000 192.080 ;
        RECT 124.180 186.620 124.510 190.470 ;
        RECT 111.940 183.470 114.750 183.955 ;
        RECT 108.000 182.790 108.260 183.130 ;
        RECT 108.515 183.110 118.395 183.470 ;
        RECT 113.210 182.790 113.470 182.800 ;
        RECT 118.640 182.790 118.900 183.130 ;
        RECT 108.000 182.530 118.900 182.790 ;
        RECT 108.000 182.190 108.260 182.530 ;
        RECT 104.570 180.560 112.450 180.610 ;
        RECT 87.420 180.300 99.340 180.560 ;
        RECT 100.670 180.300 112.450 180.560 ;
        RECT 87.420 180.250 95.300 180.300 ;
        RECT 104.570 180.250 112.450 180.300 ;
        RECT 113.210 179.000 113.470 182.530 ;
        RECT 118.640 182.190 118.900 182.530 ;
        RECT 114.230 180.560 122.110 180.610 ;
        RECT 125.760 180.560 126.020 194.560 ;
        RECT 132.940 193.750 136.520 194.040 ;
        RECT 127.890 192.780 146.850 193.580 ;
        RECT 132.710 191.770 133.600 192.440 ;
        RECT 127.890 185.490 146.850 186.290 ;
        RECT 131.270 184.010 131.680 184.550 ;
        RECT 135.780 184.010 136.170 184.610 ;
        RECT 131.270 183.600 136.170 184.010 ;
        RECT 131.270 182.980 131.680 183.600 ;
        RECT 114.230 180.300 126.150 180.560 ;
        RECT 114.230 180.250 122.110 180.300 ;
        RECT 73.730 178.740 86.660 179.000 ;
        RECT 100.540 178.740 113.470 179.000 ;
        RECT 127.890 178.200 146.850 179.000 ;
        RECT 73.730 177.620 86.660 177.880 ;
        RECT 100.540 177.620 113.470 177.880 ;
        RECT 77.760 176.320 85.640 176.370 ;
        RECT 73.860 176.060 85.640 176.320 ;
        RECT 73.860 162.060 74.120 176.060 ;
        RECT 77.760 176.010 85.640 176.060 ;
        RECT 81.190 174.090 81.450 174.430 ;
        RECT 86.400 174.090 86.660 177.620 ;
        RECT 87.420 176.320 95.300 176.370 ;
        RECT 104.570 176.320 112.450 176.370 ;
        RECT 87.420 176.060 99.340 176.320 ;
        RECT 100.670 176.060 112.450 176.320 ;
        RECT 87.420 176.010 95.300 176.060 ;
        RECT 91.830 174.090 92.090 174.430 ;
        RECT 81.190 173.830 92.090 174.090 ;
        RECT 81.190 173.490 81.450 173.830 ;
        RECT 86.400 173.820 86.660 173.830 ;
        RECT 81.705 173.150 91.585 173.510 ;
        RECT 91.830 173.490 92.090 173.830 ;
        RECT 85.130 172.665 87.940 173.150 ;
        RECT 75.370 169.640 75.710 172.360 ;
        RECT 75.370 167.590 75.700 169.640 ;
        RECT 75.370 167.240 75.710 167.590 ;
        RECT 75.880 164.540 76.600 170.850 ;
        RECT 77.080 165.680 77.800 169.640 ;
        RECT 85.140 167.590 85.860 172.665 ;
        RECT 86.000 167.240 86.340 172.360 ;
        RECT 86.730 166.150 87.070 169.990 ;
        RECT 87.220 167.570 87.940 172.665 ;
        RECT 77.540 164.960 77.800 165.680 ;
        RECT 95.270 165.350 95.990 169.620 ;
        RECT 95.270 165.300 95.940 165.350 ;
        RECT 80.690 164.960 80.950 164.970 ;
        RECT 95.270 164.960 95.530 165.300 ;
        RECT 77.540 164.700 80.950 164.960 ;
        RECT 80.690 164.540 80.950 164.700 ;
        RECT 92.280 164.700 95.530 164.960 ;
        RECT 92.280 164.540 92.540 164.700 ;
        RECT 96.470 164.540 97.190 170.860 ;
        RECT 97.370 166.150 97.700 170.000 ;
        RECT 74.840 164.180 78.720 164.540 ;
        RECT 80.690 164.180 85.570 164.540 ;
        RECT 87.660 164.180 92.540 164.540 ;
        RECT 94.340 164.180 98.220 164.540 ;
        RECT 80.690 162.060 85.570 162.110 ;
        RECT 73.860 161.800 85.570 162.060 ;
        RECT 80.690 161.750 85.570 161.800 ;
        RECT 85.770 160.810 86.030 164.180 ;
        RECT 87.200 160.810 87.460 164.180 ;
        RECT 87.660 162.060 92.540 162.110 ;
        RECT 98.950 162.060 99.210 176.060 ;
        RECT 87.660 161.800 99.210 162.060 ;
        RECT 100.670 162.060 100.930 176.060 ;
        RECT 104.570 176.010 112.450 176.060 ;
        RECT 108.000 174.090 108.260 174.430 ;
        RECT 113.210 174.090 113.470 177.620 ;
        RECT 114.230 176.320 122.110 176.370 ;
        RECT 114.230 176.060 126.150 176.320 ;
        RECT 114.230 176.010 122.110 176.060 ;
        RECT 118.640 174.090 118.900 174.430 ;
        RECT 108.000 173.830 118.900 174.090 ;
        RECT 108.000 173.490 108.260 173.830 ;
        RECT 113.210 173.820 113.470 173.830 ;
        RECT 108.515 173.150 118.395 173.510 ;
        RECT 118.640 173.490 118.900 173.830 ;
        RECT 111.940 172.665 114.750 173.150 ;
        RECT 102.180 169.640 102.520 172.360 ;
        RECT 102.180 167.590 102.510 169.640 ;
        RECT 102.180 167.240 102.520 167.590 ;
        RECT 102.690 164.540 103.410 170.850 ;
        RECT 103.890 165.680 104.610 169.640 ;
        RECT 111.950 167.590 112.670 172.665 ;
        RECT 112.810 167.240 113.150 172.360 ;
        RECT 113.540 166.150 113.880 169.990 ;
        RECT 114.030 167.570 114.750 172.665 ;
        RECT 104.350 164.960 104.610 165.680 ;
        RECT 122.080 165.350 122.800 169.620 ;
        RECT 122.080 165.300 122.750 165.350 ;
        RECT 107.500 164.960 107.760 164.970 ;
        RECT 122.080 164.960 122.340 165.300 ;
        RECT 104.350 164.700 107.760 164.960 ;
        RECT 107.500 164.540 107.760 164.700 ;
        RECT 119.090 164.700 122.340 164.960 ;
        RECT 119.090 164.540 119.350 164.700 ;
        RECT 123.280 164.540 124.000 170.860 ;
        RECT 124.180 166.150 124.510 170.000 ;
        RECT 101.650 164.180 105.530 164.540 ;
        RECT 107.500 164.180 112.380 164.540 ;
        RECT 114.470 164.180 119.350 164.540 ;
        RECT 121.150 164.180 125.030 164.540 ;
        RECT 107.500 162.060 112.380 162.110 ;
        RECT 100.670 161.800 112.380 162.060 ;
        RECT 87.660 161.750 92.540 161.800 ;
        RECT 107.500 161.750 112.380 161.800 ;
        RECT 112.580 160.810 112.840 164.180 ;
        RECT 114.010 160.810 114.270 164.180 ;
        RECT 114.470 162.060 119.350 162.110 ;
        RECT 125.760 162.060 126.020 176.060 ;
        RECT 131.250 173.600 131.700 174.200 ;
        RECT 131.250 173.180 135.360 173.600 ;
        RECT 131.250 172.630 131.700 173.180 ;
        RECT 127.890 170.910 146.850 171.710 ;
        RECT 131.240 168.820 131.670 169.930 ;
        RECT 131.240 168.380 136.930 168.820 ;
        RECT 127.890 164.020 146.850 164.420 ;
        RECT 114.470 161.800 126.020 162.060 ;
        RECT 114.470 161.750 119.350 161.800 ;
        RECT 107.490 157.800 112.370 157.850 ;
        RECT 100.660 157.540 112.370 157.800 ;
        RECT 100.660 143.540 100.920 157.540 ;
        RECT 107.490 157.490 112.370 157.540 ;
        RECT 112.570 155.420 112.830 158.790 ;
        RECT 114.000 155.420 114.260 158.790 ;
        RECT 114.460 157.800 119.340 157.850 ;
        RECT 114.460 157.540 126.010 157.800 ;
        RECT 114.460 157.490 119.340 157.540 ;
        RECT 101.640 155.060 105.520 155.420 ;
        RECT 107.490 155.060 112.370 155.420 ;
        RECT 114.460 155.060 119.340 155.420 ;
        RECT 121.140 155.060 125.020 155.420 ;
        RECT 102.170 152.010 102.510 152.360 ;
        RECT 102.170 149.960 102.500 152.010 ;
        RECT 102.170 147.240 102.510 149.960 ;
        RECT 102.680 148.750 103.400 155.060 ;
        RECT 107.490 154.900 107.750 155.060 ;
        RECT 104.340 154.640 107.750 154.900 ;
        RECT 119.080 154.900 119.340 155.060 ;
        RECT 119.080 154.640 122.330 154.900 ;
        RECT 104.340 153.920 104.600 154.640 ;
        RECT 107.490 154.630 107.750 154.640 ;
        RECT 103.880 149.960 104.600 153.920 ;
        RECT 122.070 154.300 122.330 154.640 ;
        RECT 122.070 154.250 122.740 154.300 ;
        RECT 111.940 146.935 112.660 152.010 ;
        RECT 112.800 147.240 113.140 152.360 ;
        RECT 113.530 149.610 113.870 153.450 ;
        RECT 114.020 146.935 114.740 152.030 ;
        RECT 122.070 149.980 122.790 154.250 ;
        RECT 123.270 148.740 123.990 155.060 ;
        RECT 124.170 149.600 124.500 153.450 ;
        RECT 111.930 146.450 114.740 146.935 ;
        RECT 107.990 145.770 108.250 146.110 ;
        RECT 108.505 146.090 118.385 146.450 ;
        RECT 113.200 145.770 113.460 145.780 ;
        RECT 118.630 145.770 118.890 146.110 ;
        RECT 107.990 145.510 118.890 145.770 ;
        RECT 107.990 145.170 108.250 145.510 ;
        RECT 104.560 143.540 112.440 143.590 ;
        RECT 100.660 143.280 112.440 143.540 ;
        RECT 104.560 143.230 112.440 143.280 ;
        RECT 113.200 141.980 113.460 145.510 ;
        RECT 118.630 145.170 118.890 145.510 ;
        RECT 114.220 143.540 122.100 143.590 ;
        RECT 125.750 143.540 126.010 157.540 ;
        RECT 114.220 143.280 126.140 143.540 ;
        RECT 114.220 143.230 122.100 143.280 ;
        RECT 100.530 141.720 113.460 141.980 ;
      LAYER met3 ;
        RECT 129.190 164.020 131.790 215.050 ;
        RECT 136.560 212.770 136.950 213.750 ;
        RECT 136.560 212.280 137.810 212.770 ;
        RECT 132.970 192.430 133.320 210.920 ;
        RECT 134.980 202.300 135.360 202.310 ;
        RECT 136.530 202.300 136.960 203.260 ;
        RECT 134.980 201.880 136.960 202.300 ;
        RECT 132.760 191.800 133.560 192.430 ;
        RECT 134.980 173.600 135.360 201.880 ;
        RECT 137.420 201.170 137.810 212.280 ;
        RECT 139.390 205.840 139.770 212.240 ;
        RECT 140.580 205.310 141.020 211.070 ;
        RECT 135.780 200.850 137.810 201.170 ;
        RECT 135.780 183.600 136.170 200.850 ;
        RECT 134.070 173.180 135.360 173.600 ;
        RECT 136.560 168.820 136.930 198.220 ;
        RECT 135.430 168.380 136.930 168.820 ;
        RECT 138.260 164.020 141.210 200.870 ;
        RECT 141.850 198.680 142.220 206.580 ;
        RECT 143.180 164.020 145.920 215.050 ;
  END
END tt_um_tinyflash
END LIBRARY

