magic
tech sky130A
magscale 1 2
timestamp 1762640459
<< viali >>
rect 128 802 1096 836
rect 138 -566 1106 -532
<< metal1 >>
rect 86 836 1140 872
rect 86 802 128 836
rect 1096 802 1140 836
rect 86 792 1140 802
rect 118 642 184 792
rect 264 694 646 750
rect 896 696 962 750
rect 118 264 270 642
rect 324 266 446 642
rect 264 -142 330 210
rect 394 68 446 266
rect 482 266 586 642
rect 388 64 454 68
rect 388 4 396 64
rect 448 4 454 64
rect 388 -2 454 4
rect 394 -188 446 -2
rect 112 -364 270 -188
rect 324 -364 446 -188
rect 482 -188 518 266
rect 640 264 902 642
rect 956 264 1080 642
rect 580 156 646 212
rect 580 8 586 66
rect 640 8 646 66
rect 580 -144 646 8
rect 708 -188 834 264
rect 896 64 962 212
rect 896 8 898 64
rect 960 8 962 64
rect 896 2 962 8
rect 896 -140 962 -88
rect 1024 -188 1080 264
rect 482 -364 586 -188
rect 640 -364 902 -188
rect 956 -364 1080 -188
rect 112 -506 170 -364
rect 244 -416 350 -410
rect 244 -468 260 -416
rect 332 -468 350 -416
rect 580 -464 646 -410
rect 874 -418 980 -410
rect 244 -476 350 -468
rect 874 -470 892 -418
rect 964 -470 980 -418
rect 874 -476 980 -470
rect 86 -532 1140 -506
rect 86 -566 138 -532
rect 1106 -566 1140 -532
rect 86 -586 1140 -566
<< via1 >>
rect 396 4 448 64
rect 586 8 640 66
rect 898 8 960 64
rect 260 -468 332 -416
rect 892 -470 964 -418
<< metal2 >>
rect 388 66 966 68
rect 388 64 586 66
rect 388 4 396 64
rect 448 8 586 64
rect 640 64 966 66
rect 640 8 898 64
rect 960 8 966 64
rect 448 4 966 8
rect 388 2 966 4
rect 254 -416 970 -414
rect 254 -468 260 -416
rect 332 -418 970 -416
rect 332 -468 892 -418
rect 254 -470 892 -468
rect 964 -470 970 -418
rect 254 -472 970 -470
use sky130_fd_pr__pfet_01v8_A6MZLZ  XM1
timestamp 1762640459
transform 1 0 297 0 1 453
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_MH3LLV  XM2
timestamp 1762640459
transform 1 0 297 0 1 -276
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_A6MZLZ  XM3
timestamp 1762640459
transform 1 0 613 0 1 453
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_MH3LLV  XM4
timestamp 1762640459
transform 1 0 613 0 1 -276
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_A6MZLZ  XM5
timestamp 1762640459
transform 1 0 929 0 1 453
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_MH3LLV  XM6
timestamp 1762640459
transform 1 0 929 0 1 -276
box -211 -310 211 310
<< labels >>
rlabel metal1 482 266 586 642 1 A
port 0 n
rlabel metal1 956 264 1080 642 1 B
port 1 n
rlabel metal1 264 -142 330 210 1 S
port 2 n
rlabel metal1 640 -364 902 -188 1 Y
port 3 n
rlabel metal1 86 836 1140 872 1 vdd
port 4 n
rlabel metal1 86 -586 122 -520 1 vss
port 5 n
<< end >>
