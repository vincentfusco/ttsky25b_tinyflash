* NGSPICE file created from tt_um_tinyflash_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9 B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_1p41 l=7
C0 R2 R1 0.01316f
C1 R2 B 0.87037f
C2 R1 B 0.87037f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ELBHUY B D S G
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 G D 0.11229f
C1 S D 0.27388f
C2 S G 0.11229f
C3 S B 0.59197f
C4 D B 0.59197f
C5 G B 0.75059f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_VTBKAA D S G w_n200_n1220# VSUBS
X0 S G D w_n200_n1220# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 S G 0.21915f
C1 S w_n200_n1220# 0.62529f
C2 w_n200_n1220# G 0.28692f
C3 D S 0.54671f
C4 D G 0.21915f
C5 D w_n200_n1220# 0.04108f
C6 S VSUBS 0.52213f
C7 D VSUBS 0.93676f
C8 G VSUBS 0.45532f
C9 w_n200_n1220# VSUBS 4.23183f
.ends

.subckt vbias_generation bias_n XR_bias_2/R2 XR_bias_1/R2 XR_bias_4/R1 vdd XR_bias_3/R2
+ bias_p vss
XXR_bias_1 vss XR_bias_2/R2 XR_bias_1/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_2 vss XR_bias_3/R2 XR_bias_2/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_3 vss XR_bias_4/R1 XR_bias_3/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_4 vss XR_bias_4/R1 bias_n sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXMn_bias vss bias_n vss bias_n sky130_fd_pr__nfet_01v8_lvt_ELBHUY
XXMp_bias bias_p vdd bias_p vdd vss sky130_fd_pr__pfet_01v8_lvt_VTBKAA
C0 XR_bias_3/R2 XR_bias_1/R2 0.1119f
C1 vdd XR_bias_1/R2 0.00287f
C2 XR_bias_2/R2 XR_bias_4/R1 0.1119f
C3 XR_bias_3/R2 bias_n 0.11211f
C4 XR_bias_3/R2 bias_p 0
C5 vdd bias_p 0.11094f
C6 bias_p XR_bias_1/R2 0.05695f
C7 XR_bias_3/R2 XR_bias_4/R1 0
C8 XR_bias_3/R2 XR_bias_2/R2 0
C9 XR_bias_2/R2 vdd 0.01298f
C10 XR_bias_2/R2 XR_bias_1/R2 0
C11 XR_bias_4/R1 bias_n 0
C12 XR_bias_4/R1 bias_p 0
C13 XR_bias_2/R2 bias_p 0.04272f
C14 vdd vss 5.12115f
C15 bias_p vss 1.25296f
C16 bias_n vss 2.50406f
C17 XR_bias_4/R1 vss 1.66866f
C18 XR_bias_3/R2 vss 1.56208f
C19 XR_bias_2/R2 vss 1.60214f
C20 XR_bias_1/R2 vss 0.76544f
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_JT48NU B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_5p73 l=5.73
C0 R1 R2 0.06813f
C1 R2 B 1.79077f
C2 R1 B 1.79077f
.ends

.subckt res_ladder_vref ref2 ref5 ref6 vref ref3 ref1 ref0 ref4 vss
XXR1 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR2 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR10 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR3 vss ref6 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR4 vss ref4 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR5 vss ref4 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR6 vss ref2 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR7 vss ref2 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR8 vss ref0 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR9 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
C0 ref1 ref0 0
C1 vss ref1 0.25149f
C2 vref ref6 0.16095f
C3 ref3 ref5 0.11224f
C4 vref ref5 0.11224f
C5 ref3 ref4 0
C6 ref3 vss 0.13925f
C7 ref2 ref0 0.11224f
C8 ref2 ref4 0.11224f
C9 vss vref 0.56362f
C10 vss ref2 0.13925f
C11 ref6 ref5 0
C12 ref3 ref1 0.11224f
C13 ref6 ref4 0.11224f
C14 vss ref6 0.25998f
C15 ref1 ref2 0
C16 ref4 ref5 0
C17 vss ref5 0.13925f
C18 vss ref0 0.4239f
C19 vss ref4 0.13925f
C20 ref3 ref2 0
C21 vss 0 -4.81991f
C22 ref1 0 3.26193f
C23 ref2 0 3.26193f
C24 ref3 0 3.26193f
C25 ref4 0 3.26193f
C26 ref5 0 3.26193f
C27 ref6 0 4.96136f
C28 ref0 0 4.96062f
C29 vref 0 4.20822f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MMMA4V a_n260_n698# a_100_n500# a_n158_n500# a_n100_n588#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n698# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 a_100_n500# a_n158_n500# 0.27388f
C1 a_100_n500# a_n100_n588# 0.11229f
C2 a_n100_n588# a_n158_n500# 0.11229f
C3 a_100_n500# a_n260_n698# 0.5905f
C4 a_n158_n500# a_n260_n698# 0.5905f
C5 a_n100_n588# a_n260_n698# 0.7183f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_5VNMZ8 a_n100_n897# a_100_n800# w_n296_n1019#
+ a_n158_n800# VSUBS
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n296_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
C0 a_n158_n800# a_100_n800# 0.43758f
C1 a_n158_n800# a_n100_n897# 0.17641f
C2 a_100_n800# a_n100_n897# 0.17641f
C3 a_n158_n800# w_n296_n1019# 0.51205f
C4 a_100_n800# w_n296_n1019# 0.51205f
C5 w_n296_n1019# a_n100_n897# 0.43443f
C6 a_100_n800# VSUBS 0.41369f
C7 a_n158_n800# VSUBS 0.41369f
C8 a_n100_n897# VSUBS 0.36418f
C9 w_n296_n1019# VSUBS 4.82082f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHMAL2 a_n260_n574# a_100_n400# a_n158_n400# a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n260_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
C0 a_100_n400# a_n158_n400# 0.21931f
C1 a_100_n400# a_n100_n488# 0.09092f
C2 a_n100_n488# a_n158_n400# 0.09092f
C3 a_100_n400# a_n260_n574# 0.48057f
C4 a_n158_n400# a_n260_n574# 0.48057f
C5 a_n100_n488# a_n260_n574# 0.74751f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GUWLND a_n158_n1000# a_n100_n1097# w_n296_n1219#
+ a_100_n1000# VSUBS
X0 a_100_n1000# a_n100_n1097# a_n158_n1000# w_n296_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 a_n158_n1000# a_100_n1000# 0.54671f
C1 a_n158_n1000# a_n100_n1097# 0.21915f
C2 a_100_n1000# a_n100_n1097# 0.21915f
C3 a_n158_n1000# w_n296_n1219# 0.634f
C4 a_100_n1000# w_n296_n1219# 0.634f
C5 w_n296_n1219# a_n100_n1097# 0.43443f
C6 a_100_n1000# VSUBS 0.51455f
C7 a_n158_n1000# VSUBS 0.51455f
C8 a_n100_n1097# VSUBS 0.36418f
C9 w_n296_n1219# VSUBS 5.72384f
.ends

.subckt comp_p vinp vinn vbias_p vdd tail vout latch_right out_left latch_left vss
XXMn_cs_left vss latch_right vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_out out_left vdd vdd vout vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_diode_left1 vss latch_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_AHMAL2
XXMn_cs_right1 vss latch_left vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_diode_right vss latch_right vss latch_right sky130_fd_pr__nfet_01v8_lvt_AHMAL2
Xsky130_fd_pr__pfet_01v8_lvt_5VNMZ8_0 out_left vdd vdd out_left vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_out_left vss out_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_out_right vss vout vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_tail tail vbias_p vdd vdd vss sky130_fd_pr__pfet_01v8_lvt_GUWLND
X0 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X1 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X2 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X3 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X4 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X5 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X6 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X7 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
C0 vinp out_left 0.22514f
C1 vinp vdd 4.26352f
C2 vbias_p out_left 0.84152f
C3 vinn latch_right 3.53507f
C4 vbias_p vdd 2.11961f
C5 vout vinn 0.12978f
C6 tail latch_right 8.8942f
C7 vout tail 0.00803f
C8 vinn latch_left 1.33911f
C9 vinp vbias_p 0.03011f
C10 latch_right out_left 0.1431f
C11 latch_right vdd 1.44611f
C12 tail latch_left 8.82993f
C13 vout out_left 0.6058f
C14 vout vdd 1.62919f
C15 latch_left out_left 0.73463f
C16 latch_left vdd 1.3971f
C17 vinp latch_right 0.51311f
C18 vbias_p latch_right 0.00109f
C19 tail vinn 0.82695f
C20 vout vinp 0.03655f
C21 vout vbias_p 0.14426f
C22 vinp latch_left 0.5043f
C23 vbias_p latch_left 0.00103f
C24 vinn out_left 0.08183f
C25 vinn vdd 2.30474f
C26 tail out_left 0.00652f
C27 tail vdd 2.22915f
C28 vout latch_right 0.72835f
C29 vinp vinn 1.25697f
C30 latch_left latch_right 5.15792f
C31 vinn vbias_p 0.00222f
C32 vdd out_left 2.99708f
C33 vinp tail 2.91757f
C34 vout latch_left 0.14014f
C35 tail vbias_p 0.65167f
C36 vinp vss 0.4258f
C37 vinn vss 0.50566f
C38 tail vss 1.09774f
C39 vbias_p vss 0.82905f
C40 vdd vss 43.54159f
C41 vout vss 3.2381f
C42 latch_right vss 4.74799f
C43 out_left vss 3.38408f
C44 latch_left vss 5.11722f
.ends

.subckt sky130_fd_pr__pfet_01v8_A6MZLZ B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 B G 0.24043f
C1 G D 0.02934f
C2 B D 0.14266f
C3 S G 0.02934f
C4 S B 0.14266f
C5 S D 0.32105f
C6 S VSUBS 0.09023f
C7 D VSUBS 0.09023f
C8 G VSUBS 0.11914f
C9 B VSUBS 1.5811f
.ends

.subckt sky130_fd_pr__nfet_01v8_MH3LLV B D S G
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 G D 0.02545f
C1 D S 0.16211f
C2 G S 0.02545f
C3 S B 0.1317f
C4 D B 0.1317f
C5 G B 0.34289f
.ends

.subckt tmux_2to1 Y vdd XM5/G A B S vss
XXM1 vdd vdd XM5/G S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM2 vss vss XM5/G S sky130_fd_pr__nfet_01v8_MH3LLV
XXM3 vdd A Y S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM4 vss A Y XM5/G sky130_fd_pr__nfet_01v8_MH3LLV
XXM5 vdd Y B XM5/G vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM6 vss Y B S sky130_fd_pr__nfet_01v8_MH3LLV
C0 A S 0.09932f
C1 vdd Y 0.18933f
C2 vdd XM5/G 0.17343f
C3 vdd B 0.11322f
C4 vdd S 0.27839f
C5 Y XM5/G 0.31571f
C6 Y B 0.03022f
C7 A vdd 0.05809f
C8 Y S 0.13093f
C9 B XM5/G 0.09611f
C10 S XM5/G 0.4752f
C11 A Y 0.03022f
C12 S B 0.0426f
C13 A XM5/G 0.66126f
C14 B vss 0.39578f
C15 S vss 1.22376f
C16 Y vss 0.38976f
C17 XM5/G vss 0.68597f
C18 vdd vss 4.09633f
C19 A vss 0.18036f
.ends

.subckt sky130_fd_pr__res_generic_m1_SPQYYJ R1 R2 m1_n100_n100# VSUBS
R0 R1 R2 sky130_fd_pr__res_generic_m1 w=1 l=1
C0 R2 VSUBS 0.07051f
C1 R1 VSUBS 0.07051f
C2 m1_n100_n100# VSUBS 0.10692f
.ends

.subckt inv vin vdd vout vss
XXMn vss vss vout vin sky130_fd_pr__nfet_01v8_MH3LLV
XXMp vdd vdd vout vin vss sky130_fd_pr__pfet_01v8_A6MZLZ
C0 vin vout 0.12658f
C1 vdd vin 0.13776f
C2 vdd vout 0.11998f
C3 vin vss 0.56678f
C4 vout vss 0.40687f
C5 vdd vss 1.84972f
.ends

.subckt buffer in out vdd inv_1/vin vss
Xinv_0 in vdd inv_1/vin vss inv
Xinv_1 inv_1/vin vdd out vss inv
C0 vdd inv_1/vin 0.16476f
C1 vdd in 0.01965f
C2 out vdd 0.00589f
C3 in inv_1/vin 0.01628f
C4 out inv_1/vin 0.0071f
C5 inv_1/vin vss 0.60193f
C6 out vss 0.3255f
C7 in vss 0.41789f
C8 vdd vss 3.06334f
.ends

.subckt tmux_7therm_to_3bin d0 d1 d2 d3 d4 d5 d6 q0 q1 q2 buffer_7/inv_1/vin buffer_3/inv_1/vin
+ buffer_2/out buffer_8/inv_1/vin buffer_4/inv_1/vin buffer_0/inv_1/vin buffer_6/out
+ R1/R2 buffer_9/inv_1/vin buffer_0/out buffer_5/inv_1/vin buffer_5/out buffer_1/inv_1/vin
+ tmux_2to1_0/XM5/G tmux_2to1_3/B tmux_2to1_1/XM5/G tmux_2to1_3/A tmux_2to1_2/XM5/G
+ tmux_2to1_3/XM5/G R1/R1 buffer_6/inv_1/vin buffer_2/inv_1/vin R1/m1_n100_n100# buffer_1/out
+ buffer_8/in vdd vss buffer_7/in buffer_4/out
Xtmux_2to1_1 buffer_8/in vdd tmux_2to1_1/XM5/G buffer_1/out buffer_5/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_2 tmux_2to1_3/B vdd tmux_2to1_2/XM5/G buffer_2/out buffer_6/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_3 buffer_7/in vdd tmux_2to1_3/XM5/G tmux_2to1_3/A tmux_2to1_3/B buffer_8/in
+ vss tmux_2to1
XR1 R1/R1 R1/R2 R1/m1_n100_n100# vss sky130_fd_pr__res_generic_m1_SPQYYJ
Xbuffer_0 d0 buffer_0/out vdd buffer_0/inv_1/vin vss buffer
Xbuffer_1 d1 buffer_1/out vdd buffer_1/inv_1/vin vss buffer
Xbuffer_2 d2 buffer_2/out vdd buffer_2/inv_1/vin vss buffer
Xbuffer_3 d3 R1/R2 vdd buffer_3/inv_1/vin vss buffer
Xbuffer_4 d4 buffer_4/out vdd buffer_4/inv_1/vin vss buffer
Xbuffer_5 d5 buffer_5/out vdd buffer_5/inv_1/vin vss buffer
Xbuffer_6 d6 buffer_6/out vdd buffer_6/inv_1/vin vss buffer
Xbuffer_7 buffer_7/in q0 vdd buffer_7/inv_1/vin vss buffer
Xbuffer_8 buffer_8/in q1 vdd buffer_8/inv_1/vin vss buffer
Xbuffer_9 R1/R1 q2 vdd buffer_9/inv_1/vin vss buffer
Xtmux_2to1_0 tmux_2to1_3/A vdd tmux_2to1_0/XM5/G buffer_0/out buffer_4/out R1/R1 vss
+ tmux_2to1
C0 buffer_4/inv_1/vin buffer_4/out 0.0079f
C1 buffer_4/inv_1/vin buffer_5/out 0
C2 q2 tmux_2to1_3/B 0
C3 tmux_2to1_3/A buffer_7/inv_1/vin 0
C4 buffer_0/out buffer_7/in 0
C5 buffer_4/out buffer_7/inv_1/vin 0.00238f
C6 buffer_8/in buffer_7/in 0.24628f
C7 tmux_2to1_3/A d0 0
C8 vdd buffer_5/inv_1/vin 0.32846f
C9 tmux_2to1_3/A tmux_2to1_3/B 0.0101f
C10 buffer_4/out tmux_2to1_3/B 0.27941f
C11 buffer_5/out tmux_2to1_3/B 0.16421f
C12 buffer_9/inv_1/vin buffer_8/inv_1/vin 0.00438f
C13 tmux_2to1_3/A buffer_4/out 0.60354f
C14 tmux_2to1_3/A buffer_5/out 0.00456f
C15 vdd buffer_9/inv_1/vin 0.03021f
C16 buffer_4/out buffer_5/out 1.96436f
C17 tmux_2to1_3/B q1 0
C18 tmux_2to1_0/XM5/G R1/R1 0.0674f
C19 tmux_2to1_2/XM5/G R1/R1 0.26532f
C20 buffer_2/out tmux_2to1_2/XM5/G 0.14365f
C21 vdd R1/R1 2.2016f
C22 vdd d1 0.07265f
C23 buffer_0/inv_1/vin R1/R1 0.01886f
C24 vdd buffer_2/out 0.64599f
C25 buffer_2/inv_1/vin tmux_2to1_3/B 0
C26 vdd R1/m1_n100_n100# 0.01544f
C27 buffer_7/in buffer_7/inv_1/vin 0.00796f
C28 buffer_1/out tmux_2to1_1/XM5/G 0.18587f
C29 buffer_0/out tmux_2to1_0/XM5/G 0.18135f
C30 vdd d6 0.07265f
C31 buffer_8/in buffer_8/inv_1/vin 0.01384f
C32 vdd d4 0.07265f
C33 vdd d5 0.07265f
C34 buffer_4/out R1/R2 0.00232f
C35 buffer_5/out R1/R2 0.01212f
C36 buffer_7/in tmux_2to1_3/B 0.20877f
C37 buffer_0/out vdd 0.83616f
C38 buffer_0/out buffer_0/inv_1/vin 0.00873f
C39 tmux_2to1_3/XM5/G R1/R1 0
C40 buffer_8/in vdd 0.52301f
C41 tmux_2to1_3/A buffer_7/in 0.38438f
C42 buffer_7/in buffer_4/out 0.04488f
C43 buffer_7/in buffer_5/out 0.00264f
C44 buffer_5/inv_1/vin buffer_6/out 0
C45 buffer_8/in tmux_2to1_3/XM5/G 0.34642f
C46 buffer_2/inv_1/vin buffer_1/inv_1/vin 0.00438f
C47 buffer_7/in q1 0
C48 buffer_4/inv_1/vin vdd 0.32846f
C49 tmux_2to1_3/A q0 0
C50 buffer_8/inv_1/vin buffer_7/inv_1/vin 0.00435f
C51 buffer_9/inv_1/vin buffer_6/out 0.00222f
C52 buffer_8/inv_1/vin tmux_2to1_3/B 0.00974f
C53 d0 tmux_2to1_0/XM5/G 0
C54 vdd buffer_7/inv_1/vin 0.02382f
C55 tmux_2to1_2/XM5/G tmux_2to1_3/B 0.03416f
C56 buffer_3/inv_1/vin R1/R1 0.00894f
C57 vdd d0 0.0683f
C58 vdd tmux_2to1_3/B 1.44834f
C59 buffer_6/out R1/R1 0.20693f
C60 vdd q2 0.01294f
C61 tmux_2to1_3/A tmux_2to1_0/XM5/G 0.08101f
C62 buffer_2/out buffer_6/out 0.01539f
C63 buffer_3/inv_1/vin R1/m1_n100_n100# 0.00103f
C64 buffer_5/out buffer_8/inv_1/vin 0
C65 R1/m1_n100_n100# buffer_6/out 0
C66 buffer_4/out tmux_2to1_0/XM5/G 0.02654f
C67 buffer_4/out tmux_2to1_2/XM5/G 0.07683f
C68 buffer_5/out tmux_2to1_2/XM5/G 0.09828f
C69 d6 buffer_6/out 0.00132f
C70 tmux_2to1_3/A vdd 0.31099f
C71 tmux_2to1_3/A buffer_0/inv_1/vin 0
C72 vdd buffer_4/out 1.78677f
C73 vdd buffer_5/out 1.96257f
C74 tmux_2to1_3/XM5/G tmux_2to1_3/B 0.0457f
C75 buffer_1/out R1/R1 0.22519f
C76 buffer_1/out d1 0.00148f
C77 vdd d3 0.07265f
C78 q0 buffer_7/in 0
C79 tmux_2to1_3/A tmux_2to1_3/XM5/G 0.04146f
C80 vdd q1 0.01294f
C81 buffer_4/out tmux_2to1_3/XM5/G 0.04713f
C82 buffer_5/out tmux_2to1_3/XM5/G 0.01262f
C83 tmux_2to1_1/XM5/G R1/R1 0.13419f
C84 vdd buffer_1/inv_1/vin 0.32649f
C85 buffer_1/inv_1/vin buffer_0/inv_1/vin 0.00435f
C86 buffer_8/in buffer_1/out 0.06403f
C87 vdd R1/R2 0.32828f
C88 vdd buffer_2/inv_1/vin 0.32649f
C89 buffer_7/in buffer_8/inv_1/vin 0
C90 buffer_7/in tmux_2to1_0/XM5/G 0.00597f
C91 R1/R1 d2 0.00119f
C92 d1 d2 0.00438f
C93 buffer_4/inv_1/vin buffer_3/inv_1/vin 0.00438f
C94 buffer_4/inv_1/vin buffer_6/out 0
C95 buffer_2/out d2 0
C96 buffer_8/in tmux_2to1_1/XM5/G 0.12457f
C97 vdd buffer_6/inv_1/vin 0.32835f
C98 vdd buffer_7/in 0.23539f
C99 buffer_6/out tmux_2to1_3/B 0.18281f
C100 buffer_7/in tmux_2to1_3/XM5/G 0.01403f
C101 buffer_4/out buffer_3/inv_1/vin 0
C102 buffer_3/inv_1/vin buffer_5/out 0
C103 q0 vdd 0.01294f
C104 buffer_4/out buffer_6/out 1.41966f
C105 buffer_5/out buffer_6/out 0.48773f
C106 buffer_1/out tmux_2to1_3/B 0
C107 tmux_2to1_3/A buffer_1/out 0
C108 buffer_9/inv_1/vin R1/R1 0.00349f
C109 vdd buffer_8/inv_1/vin 0.02538f
C110 vdd tmux_2to1_0/XM5/G 0.05854f
C111 vdd tmux_2to1_2/XM5/G 0.05427f
C112 tmux_2to1_1/XM5/G tmux_2to1_3/B 0
C113 buffer_1/out buffer_4/out 0.00456f
C114 buffer_1/out buffer_5/out 0.05669f
C115 tmux_2to1_0/XM5/G buffer_0/inv_1/vin 0
C116 R1/R2 buffer_6/out 0.00154f
C117 vdd buffer_0/inv_1/vin 0.32203f
C118 tmux_2to1_3/A tmux_2to1_1/XM5/G 0
C119 buffer_3/inv_1/vin buffer_2/inv_1/vin 0.00435f
C120 d2 tmux_2to1_3/B 0
C121 d1 R1/R1 0
C122 buffer_4/out tmux_2to1_1/XM5/G 0.02598f
C123 buffer_5/out tmux_2to1_1/XM5/G 0.02579f
C124 buffer_2/out R1/R1 0.2789f
C125 R1/m1_n100_n100# R1/R1 0.04565f
C126 buffer_6/inv_1/vin buffer_6/out 0.00786f
C127 buffer_1/out buffer_1/inv_1/vin 0.0086f
C128 vdd tmux_2to1_3/XM5/G 0.0495f
C129 buffer_0/out R1/R1 0.11396f
C130 buffer_4/inv_1/vin buffer_5/inv_1/vin 0.00435f
C131 buffer_8/in R1/R1 0.07792f
C132 buffer_8/in d1 0
C133 d5 d6 0.00438f
C134 d4 d5 0.00435f
C135 d3 d2 0.00435f
C136 buffer_1/out buffer_7/in 0
C137 buffer_7/in tmux_2to1_1/XM5/G 0
C138 buffer_5/out buffer_5/inv_1/vin 0.00827f
C139 buffer_9/inv_1/vin tmux_2to1_3/B 0.00176f
C140 tmux_2to1_2/XM5/G buffer_6/out 0.02333f
C141 vdd buffer_3/inv_1/vin 0.32836f
C142 vdd buffer_6/out 3.00774f
C143 d0 d1 0.00435f
C144 d0 R1/R1 0
C145 R1/R1 tmux_2to1_3/B 0.24354f
C146 q2 R1/R1 0
C147 buffer_2/out tmux_2to1_3/B 0.04026f
C148 tmux_2to1_3/A R1/R1 0.0222f
C149 buffer_4/out R1/R1 0.26729f
C150 buffer_1/out vdd 0.83708f
C151 buffer_5/out R1/R1 0.55887f
C152 buffer_0/out d0 0.0015f
C153 buffer_4/out buffer_2/out 0.0018f
C154 buffer_5/out buffer_2/out 0.05213f
C155 buffer_8/in tmux_2to1_3/B 0.28179f
C156 buffer_4/out R1/m1_n100_n100# 0.00131f
C157 buffer_5/out R1/m1_n100_n100# 0.01185f
C158 tmux_2to1_0/XM5/G tmux_2to1_1/XM5/G 0.00433f
C159 tmux_2to1_2/XM5/G tmux_2to1_1/XM5/G 0.00433f
C160 buffer_6/inv_1/vin buffer_5/inv_1/vin 0.00438f
C161 d4 buffer_4/out 0.00133f
C162 d5 buffer_5/out 0.00133f
C163 tmux_2to1_3/A buffer_0/out 0.05826f
C164 d3 R1/R1 0
C165 vdd tmux_2to1_1/XM5/G 0.04059f
C166 tmux_2to1_3/A buffer_8/in 0.1382f
C167 buffer_0/out buffer_4/out 0.0414f
C168 buffer_8/in buffer_4/out 0.18314f
C169 buffer_1/out tmux_2to1_3/XM5/G 0
C170 buffer_8/in buffer_5/out 0.33947f
C171 buffer_1/inv_1/vin R1/R1 0.02062f
C172 d4 d3 0.00438f
C173 R1/R2 R1/R1 0.03366f
C174 vdd d2 0.07265f
C175 R1/R2 R1/m1_n100_n100# 0.0386f
C176 buffer_2/inv_1/vin R1/R1 0.02182f
C177 buffer_2/inv_1/vin buffer_2/out 0.00356f
C178 buffer_8/in q1 0
C179 buffer_8/in buffer_1/inv_1/vin 0
C180 buffer_7/in R1/R1 0.00295f
C181 buffer_3/inv_1/vin buffer_6/out 0
C182 tmux_2to1_3/A vss 0.7137f
C183 tmux_2to1_0/XM5/G vss 0.55203f
C184 buffer_9/inv_1/vin vss 0.83718f
C185 q2 vss 0.40182f
C186 buffer_8/inv_1/vin vss 0.83586f
C187 q1 vss 0.40182f
C188 buffer_7/inv_1/vin vss 0.83588f
C189 q0 vss 0.40182f
C190 buffer_6/inv_1/vin vss 0.54713f
C191 buffer_6/out vss 1.08087f
C192 d6 vss 0.42023f
C193 buffer_5/inv_1/vin vss 0.54811f
C194 buffer_5/out vss 1.1426f
C195 d5 vss 0.41693f
C196 vdd vss 81.61826f
C197 buffer_4/inv_1/vin vss 0.54811f
C198 buffer_4/out vss 1.13891f
C199 d4 vss 0.41693f
C200 buffer_3/inv_1/vin vss 0.54811f
C201 R1/R2 vss 0.24596f
C202 d3 vss 0.41694f
C203 buffer_2/inv_1/vin vss 0.55981f
C204 buffer_2/out vss 0.38944f
C205 d2 vss 0.41693f
C206 buffer_1/inv_1/vin vss 0.55981f
C207 buffer_1/out vss 0.403f
C208 d1 vss 0.41693f
C209 buffer_0/inv_1/vin vss 0.55981f
C210 buffer_0/out vss 0.40723f
C211 d0 vss 0.42457f
C212 R1/m1_n100_n100# vss 0.11104f
C213 buffer_8/in vss 1.94693f
C214 buffer_7/in vss 1.30882f
C215 tmux_2to1_3/XM5/G vss 0.55181f
C216 R1/R1 vss 4.97015f
C217 tmux_2to1_3/B vss 1.00035f
C218 tmux_2to1_2/XM5/G vss 0.54992f
C219 tmux_2to1_1/XM5/G vss 0.55178f
.ends

.subckt flashADC_3bit dout0 dout1 dout2 tmux_7therm_to_3bin_0/buffer_1/out vbias_generation_0/bias_n
+ tmux_7therm_to_3bin_0/buffer_6/inv_1/vin tmux_7therm_to_3bin_0/buffer_2/inv_1/vin
+ comp_p_3/latch_left comp_p_5/tail tmux_7therm_to_3bin_0/buffer_8/in comp_p_2/tail
+ comp_p_4/latch_left tmux_7therm_to_3bin_0/buffer_7/in comp_p_5/latch_left vbias_generation_0/XR_bias_2/R2
+ tmux_7therm_to_3bin_0/R1/m1_n100_n100# tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_2/out tmux_7therm_to_3bin_0/buffer_3/inv_1/vin comp_p_6/latch_left
+ comp_p_1/out_left comp_p_6/tail comp_p_0/latch_right comp_p_1/latch_right comp_p_2/latch_right
+ comp_p_3/latch_right comp_p_3/tail comp_p_4/latch_right comp_p_5/latch_right tmux_7therm_to_3bin_0/buffer_8/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_6/out comp_p_4/out_left comp_p_4/vinn comp_p_6/latch_right
+ comp_p_0/tail tmux_7therm_to_3bin_0/buffer_4/inv_1/vin tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ tmux_7therm_to_3bin_0/R1/R2 comp_p_2/latch_left vbias_generation_0/XR_bias_4/R1
+ tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G d1 comp_p_3/vinn tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G
+ comp_p_2/out_left tmux_7therm_to_3bin_0/buffer_0/out comp_p_0/out_left tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G
+ tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G comp_p_6/vinn tmux_7therm_to_3bin_0/buffer_5/out
+ d2 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin comp_p_4/tail tmux_7therm_to_3bin_0/R1/R1
+ comp_p_0/latch_left tmux_7therm_to_3bin_0/buffer_5/inv_1/vin tmux_7therm_to_3bin_0/buffer_1/inv_1/vin
+ d4 comp_p_5/vinn tmux_7therm_to_3bin_0/tmux_2to1_3/B comp_p_1/tail comp_p_0/vinn
+ vin comp_p_6/out_left tmux_7therm_to_3bin_0/tmux_2to1_3/A comp_p_1/latch_left vdd
+ tmux_7therm_to_3bin_0/buffer_4/out d5 d3 d0 comp_p_1/vinn comp_p_2/vinn vref comp_p_5/out_left
+ vbias_generation_0/XR_bias_3/R2 d6 vss comp_p_3/out_left comp_p_6/vbias_p
Xvbias_generation_0 vbias_generation_0/bias_n vbias_generation_0/XR_bias_2/R2 comp_p_6/vbias_p
+ vbias_generation_0/XR_bias_4/R1 vdd vbias_generation_0/XR_bias_3/R2 comp_p_6/vbias_p
+ vss vbias_generation
Xres_ladder_vref_0 comp_p_2/vinn comp_p_5/vinn comp_p_6/vinn vref comp_p_3/vinn comp_p_0/vinn
+ comp_p_1/vinn comp_p_4/vinn vss res_ladder_vref
Xcomp_p_1 vin comp_p_1/vinn comp_p_6/vbias_p vdd comp_p_1/tail d0 comp_p_1/latch_right
+ comp_p_1/out_left comp_p_1/latch_left vss comp_p
Xcomp_p_0 vin comp_p_0/vinn comp_p_6/vbias_p vdd comp_p_0/tail d1 comp_p_0/latch_right
+ comp_p_0/out_left comp_p_0/latch_left vss comp_p
Xcomp_p_2 vin comp_p_2/vinn comp_p_6/vbias_p vdd comp_p_2/tail d2 comp_p_2/latch_right
+ comp_p_2/out_left comp_p_2/latch_left vss comp_p
Xcomp_p_3 vin comp_p_3/vinn comp_p_6/vbias_p vdd comp_p_3/tail d3 comp_p_3/latch_right
+ comp_p_3/out_left comp_p_3/latch_left vss comp_p
Xcomp_p_4 vin comp_p_4/vinn comp_p_6/vbias_p vdd comp_p_4/tail d4 comp_p_4/latch_right
+ comp_p_4/out_left comp_p_4/latch_left vss comp_p
Xcomp_p_5 vin comp_p_5/vinn comp_p_6/vbias_p vdd comp_p_5/tail d5 comp_p_5/latch_right
+ comp_p_5/out_left comp_p_5/latch_left vss comp_p
Xcomp_p_6 vin comp_p_6/vinn comp_p_6/vbias_p vdd comp_p_6/tail d6 comp_p_6/latch_right
+ comp_p_6/out_left comp_p_6/latch_left vss comp_p
Xtmux_7therm_to_3bin_0 d0 d1 d2 d3 d4 d5 d6 dout0 dout1 dout2 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_3/inv_1/vin tmux_7therm_to_3bin_0/buffer_2/out tmux_7therm_to_3bin_0/buffer_8/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_4/inv_1/vin tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_6/out tmux_7therm_to_3bin_0/R1/R2 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_0/out tmux_7therm_to_3bin_0/buffer_5/inv_1/vin tmux_7therm_to_3bin_0/buffer_5/out
+ tmux_7therm_to_3bin_0/buffer_1/inv_1/vin tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G
+ tmux_7therm_to_3bin_0/tmux_2to1_3/B tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G tmux_7therm_to_3bin_0/tmux_2to1_3/A
+ tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G
+ tmux_7therm_to_3bin_0/R1/R1 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin tmux_7therm_to_3bin_0/buffer_2/inv_1/vin
+ tmux_7therm_to_3bin_0/R1/m1_n100_n100# tmux_7therm_to_3bin_0/buffer_1/out tmux_7therm_to_3bin_0/buffer_8/in
+ vdd vss tmux_7therm_to_3bin_0/buffer_7/in tmux_7therm_to_3bin_0/buffer_4/out tmux_7therm_to_3bin
C0 d4 d2 0.04942f
C1 comp_p_4/vinn vdd 0.03662f
C2 comp_p_4/latch_left vin 0.00664f
C3 d5 comp_p_1/out_left 0
C4 vbias_generation_0/bias_n comp_p_6/latch_right 0
C5 d4 comp_p_6/vbias_p 0.37293f
C6 d4 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C7 comp_p_1/vinn comp_p_0/vinn 0.94729f
C8 comp_p_1/vinn comp_p_1/out_left 0.19389f
C9 d2 comp_p_3/latch_right 0.09517f
C10 tmux_7therm_to_3bin_0/buffer_6/out d6 0
C11 comp_p_6/vbias_p comp_p_0/latch_left 0.37827f
C12 d0 comp_p_1/out_left -0
C13 d3 vin 0.00158f
C14 d5 comp_p_5/out_left 0
C15 d4 tmux_7therm_to_3bin_0/buffer_2/out 0
C16 comp_p_5/latch_right comp_p_6/latch_right 0.00925f
C17 d4 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin 0.00318f
C18 comp_p_1/latch_left d2 0
C19 vbias_generation_0/bias_n comp_p_6/out_left 0.00925f
C20 vdd comp_p_6/latch_right 1.95544f
C21 comp_p_5/tail d6 0
C22 d5 d2 0.04508f
C23 d1 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0.00173f
C24 d6 comp_p_5/latch_left 0.00183f
C25 comp_p_2/vinn vdd 0.04727f
C26 d6 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C27 vdd comp_p_2/out_left 0.02487f
C28 comp_p_0/latch_left comp_p_2/latch_left 0.01494f
C29 d5 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C30 d5 comp_p_6/vbias_p 0
C31 d2 comp_p_1/vinn 0.00152f
C32 comp_p_3/vinn comp_p_3/latch_left 0.00666f
C33 comp_p_6/vbias_p comp_p_1/vinn 0.38594f
C34 d0 d2 0.03281f
C35 comp_p_4/latch_right comp_p_5/out_left 0
C36 comp_p_6/vbias_p vbias_generation_0/XR_bias_4/R1 0.02724f
C37 d4 comp_p_6/latch_left 0.06068f
C38 vdd comp_p_0/vinn 0.01961f
C39 d0 comp_p_6/vbias_p 0.00465f
C40 d0 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0.00746f
C41 vdd comp_p_6/out_left 1.67021f
C42 vdd comp_p_1/out_left 1.79183f
C43 d5 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin 0
C44 comp_p_5/vinn vin 0.66275f
C45 d4 comp_p_3/latch_right 0.00133f
C46 vbias_generation_0/bias_n comp_p_6/vbias_p 0
C47 comp_p_4/latch_right comp_p_6/vbias_p 0.40389f
C48 d3 comp_p_1/tail 0
C49 tmux_7therm_to_3bin_0/R1/R1 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C50 comp_p_2/latch_right comp_p_1/vinn 0.00771f
C51 comp_p_1/vinn comp_p_2/latch_left 0.01672f
C52 d4 comp_p_1/latch_left 0
C53 comp_p_6/vinn comp_p_4/out_left 0.04948f
C54 comp_p_5/out_left vdd 1.8042f
C55 vbias_generation_0/XR_bias_3/R2 vin 0.08368f
C56 d4 d5 4.51321f
C57 d1 comp_p_3/vinn 0
C58 d6 comp_p_3/vinn 0
C59 comp_p_4/vinn comp_p_4/out_left 0.02516f
C60 d1 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0.00482f
C61 d6 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C62 d2 vdd 1.1602f
C63 d3 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0.00238f
C64 d4 comp_p_1/vinn 0
C65 comp_p_6/vbias_p vdd 12.39904f
C66 vdd tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0.00196f
C67 d5 comp_p_3/latch_right 0.00185f
C68 d4 d0 0.03391f
C69 comp_p_4/vinn comp_p_3/vinn 0
C70 comp_p_1/vinn comp_p_0/latch_left 0.15776f
C71 d4 vbias_generation_0/bias_n 0.00802f
C72 d4 comp_p_4/latch_right 0
C73 comp_p_1/latch_left d5 0
C74 vbias_generation_0/XR_bias_2/R2 vin 0.50675f
C75 vbias_generation_0/bias_n comp_p_6/latch_left 0.01259f
C76 comp_p_2/latch_right vdd 0.00592f
C77 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vdd 0.00104f
C78 vdd comp_p_2/latch_left 0
C79 d1 tmux_7therm_to_3bin_0/buffer_0/out 0
C80 comp_p_1/latch_left comp_p_1/vinn 0.0067f
C81 comp_p_1/latch_right d1 0.09536f
C82 tmux_7therm_to_3bin_0/buffer_0/out d6 0
C83 comp_p_1/latch_right d6 0.00271f
C84 vref vdd 0
C85 comp_p_2/out_left comp_p_4/out_left 0.01584f
C86 d5 comp_p_1/vinn 0
C87 d4 comp_p_5/latch_right 0.06539f
C88 d5 d0 0.04762f
C89 d6 comp_p_3/out_left 0
C90 d6 tmux_7therm_to_3bin_0/buffer_4/out 0
C91 comp_p_2/vinn comp_p_3/vinn 0.31389f
C92 comp_p_3/vinn comp_p_2/out_left 0.01462f
C93 d4 vdd 1.46229f
C94 d2 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0.00483f
C95 comp_p_6/latch_left vdd 2.04557f
C96 comp_p_0/latch_left vdd 0
C97 comp_p_2/vinn comp_p_2/tail 0
C98 comp_p_3/latch_right vdd 1.95698f
C99 vin comp_p_0/latch_right 0.21598f
C100 d1 vin 0.63586f
C101 d6 vin 0.01178f
C102 comp_p_3/vinn comp_p_0/vinn 0.53686f
C103 comp_p_4/latch_right vbias_generation_0/XR_bias_4/R1 0
C104 comp_p_6/vinn vin 1.01745f
C105 comp_p_1/latch_left vdd 2.04615f
C106 d4 tmux_7therm_to_3bin_0/buffer_6/out 0.013f
C107 comp_p_4/vinn vin 0.52728f
C108 comp_p_4/latch_right vbias_generation_0/bias_n 0
C109 d5 vdd 2.33637f
C110 comp_p_5/vinn comp_p_4/tail 0.10856f
C111 vbias_generation_0/XR_bias_3/R2 comp_p_6/tail 0
C112 comp_p_1/vinn vdd 1.45687f
C113 comp_p_6/vbias_p comp_p_4/out_left 0.69034f
C114 comp_p_2/vinn comp_p_3/out_left 0
C115 d4 comp_p_5/tail 0.00264f
C116 comp_p_3/tail d6 0
C117 d0 vdd 2.71992f
C118 d4 comp_p_5/latch_left 0.06545f
C119 d4 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C120 d2 comp_p_3/vinn 0.24742f
C121 comp_p_6/latch_left comp_p_5/latch_left 0.00925f
C122 d2 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0.00171f
C123 comp_p_6/vbias_p comp_p_3/vinn 0.38072f
C124 d1 comp_p_1/tail 0.00457f
C125 d6 comp_p_1/tail 0
C126 vbias_generation_0/bias_n vdd 0.00188f
C127 comp_p_4/latch_right vdd 0.00589f
C128 comp_p_2/vinn vin 0.52215f
C129 d2 comp_p_2/tail -0.00224f
C130 vin comp_p_2/out_left 0.0842f
C131 comp_p_6/vbias_p comp_p_2/tail 0.31443f
C132 comp_p_2/latch_right comp_p_3/vinn 0.17593f
C133 comp_p_3/vinn comp_p_2/latch_left 0.15548f
C134 d4 tmux_7therm_to_3bin_0/buffer_5/out 0.01353f
C135 comp_p_5/latch_right vdd 1.9557f
C136 d6 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C137 d5 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C138 vin comp_p_0/vinn 0.81463f
C139 tmux_7therm_to_3bin_0/buffer_0/out d2 0
C140 vin comp_p_6/out_left 0.06197f
C141 comp_p_1/latch_right d2 0.00123f
C142 vin comp_p_1/out_left 0.07139f
C143 comp_p_3/out_left comp_p_5/out_left 0.01584f
C144 d4 comp_p_3/vinn 0
C145 d2 comp_p_3/out_left 0.67197f
C146 comp_p_5/vinn comp_p_4/latch_left 0.16266f
C147 d4 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C148 comp_p_6/vbias_p comp_p_3/out_left -0.06014f
C149 comp_p_5/out_left vin 0.06043f
C150 comp_p_4/latch_right comp_p_5/latch_left 0.02598f
C151 comp_p_3/vinn comp_p_3/latch_right 0.00805f
C152 d5 tmux_7therm_to_3bin_0/buffer_5/out 0
C153 d3 tmux_7therm_to_3bin_0/R1/R2 0
C154 d2 vin 0.72189f
C155 comp_p_6/vbias_p vin 1.44148f
C156 comp_p_2/latch_right comp_p_3/out_left 0
C157 d4 tmux_7therm_to_3bin_0/buffer_0/out 0
C158 comp_p_4/out_left vbias_generation_0/XR_bias_4/R1 0
C159 d5 comp_p_3/vinn 0
C160 d4 comp_p_1/latch_right 0
C161 comp_p_5/tail vdd 0.35567f
C162 d5 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C163 comp_p_5/latch_left vdd 2.0461f
C164 comp_p_1/vinn comp_p_3/vinn 0.03321f
C165 comp_p_2/latch_right vin 0.21614f
C166 vin comp_p_2/latch_left 0.00664f
C167 d4 comp_p_3/out_left 0
C168 comp_p_1/latch_right comp_p_3/latch_right 0.00925f
C169 d4 tmux_7therm_to_3bin_0/buffer_4/out 0
C170 vin vref 0.03789f
C171 comp_p_3/tail d2 0.00272f
C172 d0 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C173 d2 comp_p_1/tail 0
C174 d4 vin 0.72855f
C175 d5 tmux_7therm_to_3bin_0/buffer_0/out 0
C176 d5 comp_p_1/latch_right 0.0019f
C177 vin comp_p_6/latch_left 0.00266f
C178 vdd comp_p_4/out_left 0.02489f
C179 d1 comp_p_0/tail -0.00224f
C180 comp_p_1/latch_right comp_p_1/vinn 0.00799f
C181 d3 comp_p_3/latch_left 0
C182 vin comp_p_0/latch_left 0.00334f
C183 d0 tmux_7therm_to_3bin_0/buffer_0/out 0
C184 d5 comp_p_3/out_left 0.02324f
C185 d5 tmux_7therm_to_3bin_0/buffer_4/out 0
C186 vdd tmux_7therm_to_3bin_0/buffer_8/in 0
C187 comp_p_3/vinn vdd 1.48772f
C188 d3 tmux_7therm_to_3bin_0/R1/R1 0
C189 d3 tmux_7therm_to_3bin_0/buffer_1/out 0
C190 comp_p_0/out_left comp_p_2/out_left 0.09264f
C191 vdd tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C192 comp_p_6/vinn comp_p_4/latch_left 0.00606f
C193 d4 comp_p_3/tail 0
C194 d5 vin 0.0056f
C195 comp_p_2/tail vdd 0.00168f
C196 comp_p_4/vinn comp_p_4/latch_left 0.00288f
C197 comp_p_0/out_left comp_p_0/vinn 0.02276f
C198 comp_p_1/vinn vin 0.97735f
C199 d4 comp_p_1/tail 0
C200 vin vbias_generation_0/XR_bias_4/R1 0.00472f
C201 d3 d1 0.11517f
C202 d3 d6 0.07956f
C203 comp_p_5/out_left comp_p_4/tail 0
C204 tmux_7therm_to_3bin_0/buffer_0/out vdd 0
C205 comp_p_1/latch_right vdd 1.96641f
C206 vbias_generation_0/bias_n vin 0.0214f
C207 comp_p_4/latch_right vin 0.21628f
C208 dout1 dout0 -0
C209 d4 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C210 d5 comp_p_3/tail 0
C211 comp_p_3/out_left vdd 1.79594f
C212 comp_p_6/vbias_p comp_p_4/tail 0.31443f
C213 tmux_7therm_to_3bin_0/buffer_4/out vdd 0.00846f
C214 d5 comp_p_1/tail 0
C215 comp_p_0/tail comp_p_1/out_left 0
C216 comp_p_0/out_left comp_p_6/vbias_p 0.68459f
C217 comp_p_5/vinn d6 0.00513f
C218 vin vdd 9.78527f
C219 comp_p_5/vinn comp_p_6/vinn 0.03037f
C220 d4 comp_p_6/tail 0.00252f
C221 d5 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C222 comp_p_4/vinn comp_p_5/vinn 0.32186f
C223 comp_p_0/out_left comp_p_2/latch_left 0.01472f
C224 vbias_generation_0/XR_bias_3/R2 comp_p_6/vinn 0.06411f
C225 d4 comp_p_4/tail -0.00224f
C226 d3 comp_p_1/out_left 0
C227 comp_p_6/vbias_p comp_p_0/tail 0.31443f
C228 comp_p_3/tail vdd 0.35691f
C229 tmux_7therm_to_3bin_0/buffer_1/out tmux_7therm_to_3bin_0/R1/R1 0
C230 vdd comp_p_1/tail 0.35563f
C231 comp_p_2/tail comp_p_3/vinn 0.14685f
C232 comp_p_6/vbias_p comp_p_4/latch_left 0.37827f
C233 comp_p_5/tail vin 0.00233f
C234 d1 comp_p_3/latch_left 0
C235 d3 comp_p_5/out_left 0.02309f
C236 d6 comp_p_3/latch_left 0
C237 comp_p_6/vinn vbias_generation_0/XR_bias_2/R2 0.00358f
C238 d3 d2 2.50136f
C239 d1 tmux_7therm_to_3bin_0/buffer_1/out 0.01311f
C240 d1 tmux_7therm_to_3bin_0/R1/R1 0.00785f
C241 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin vdd 0
C242 d3 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C243 d3 comp_p_6/vbias_p 0
C244 d6 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0
C245 d6 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0.00531f
C246 comp_p_0/out_left comp_p_1/vinn 0.04644f
C247 comp_p_3/out_left comp_p_3/vinn 0.20126f
C248 vbias_generation_0/XR_bias_3/R2 comp_p_6/out_left 0.00563f
C249 d1 comp_p_0/latch_right 0
C250 vin comp_p_4/out_left 0.0859f
C251 d3 tmux_7therm_to_3bin_0/buffer_2/out 0
C252 d1 d6 0.09f
C253 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G d0 0
C254 d3 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin 0
C255 comp_p_5/vinn comp_p_5/out_left 0.19629f
C256 comp_p_2/tail comp_p_3/out_left 0
C257 comp_p_6/tail vdd 0.3539f
C258 comp_p_3/vinn vin 0.65736f
C259 comp_p_5/vinn comp_p_6/vbias_p 0.407f
C260 d4 d3 2.88908f
C261 tmux_7therm_to_3bin_0/buffer_7/in vdd 0.0027f
C262 vdd comp_p_4/tail 0.00166f
C263 comp_p_2/tail vin 0.0104f
C264 comp_p_1/vinn comp_p_0/tail 0.10698f
C265 d3 comp_p_3/latch_right 0.0057f
C266 comp_p_0/out_left vdd 0.01217f
C267 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G vdd 0.00166f
C268 d3 tmux_7therm_to_3bin_0/R1/m1_n100_n100# 0
C269 comp_p_4/latch_left vbias_generation_0/XR_bias_4/R1 0
C270 comp_p_1/latch_left d3 0
C271 comp_p_6/vinn comp_p_6/latch_right 0.00296f
C272 d5 d3 0.16529f
C273 comp_p_3/out_left vin 0.05071f
C274 vbias_generation_0/bias_n comp_p_4/latch_left 0
C275 d4 comp_p_5/vinn 0.25734f
C276 d3 comp_p_1/vinn 0
C277 tmux_7therm_to_3bin_0/tmux_2to1_3/A d0 0
C278 d2 comp_p_3/latch_left 0.09614f
C279 comp_p_0/latch_right comp_p_0/vinn 0.00236f
C280 d1 comp_p_0/vinn -0
C281 comp_p_0/latch_right comp_p_1/out_left 0
C282 d1 comp_p_1/out_left 0.67001f
C283 d6 comp_p_1/out_left 0
C284 d3 d0 0.03225f
C285 comp_p_6/vbias_p vbias_generation_0/XR_bias_2/R2 0.02749f
C286 vdd comp_p_0/tail 0.00166f
C287 comp_p_6/vinn comp_p_6/out_left 0.14972f
C288 d2 tmux_7therm_to_3bin_0/R1/R1 0.00763f
C289 d2 tmux_7therm_to_3bin_0/buffer_1/out 0
C290 comp_p_4/latch_left vdd 0
C291 d6 comp_p_5/out_left 0
C292 comp_p_2/latch_right comp_p_3/latch_left 0.02598f
C293 comp_p_2/vinn comp_p_2/out_left 0.0232f
C294 d1 d2 3.44306f
C295 d2 comp_p_0/latch_right 0.01472f
C296 d2 d6 0.05303f
C297 tmux_7therm_to_3bin_0/tmux_2to1_3/A vdd 0.00153f
C298 comp_p_4/vinn comp_p_5/out_left 0
C299 d1 comp_p_6/vbias_p 0.37529f
C300 d1 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0.00131f
C301 comp_p_6/vbias_p comp_p_0/latch_right 0.40389f
C302 d6 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C303 d3 vdd 2.3721f
C304 comp_p_3/tail vin 0.00233f
C305 comp_p_6/vinn comp_p_6/vbias_p 0.31983f
C306 d4 comp_p_3/latch_left 0
C307 comp_p_2/vinn comp_p_0/vinn 0.02754f
C308 comp_p_2/out_left comp_p_0/vinn 0.0271f
C309 comp_p_4/latch_right comp_p_5/vinn 0.20935f
C310 vin comp_p_1/tail 0.00233f
C311 comp_p_4/vinn comp_p_6/vbias_p 0.12306f
C312 tmux_7therm_to_3bin_0/buffer_2/out d1 0.00551f
C313 d1 comp_p_2/latch_right 0.01472f
C314 comp_p_2/latch_right comp_p_0/latch_right 0.01494f
C315 d4 tmux_7therm_to_3bin_0/R1/R1 0
C316 d4 tmux_7therm_to_3bin_0/buffer_1/out 0
C317 d6 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin 0
C318 d4 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.00384f
C319 comp_p_6/vinn vref 0.00148f
C320 comp_p_1/out_left comp_p_0/vinn 0
C321 d4 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0.00248f
C322 comp_p_1/latch_left comp_p_3/latch_left 0.00925f
C323 comp_p_5/vinn comp_p_5/latch_right 0.00802f
C324 d5 comp_p_3/latch_left 0
C325 d4 d1 0.33457f
C326 comp_p_5/vinn vdd 1.45079f
C327 d4 d6 0.79887f
C328 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vdd 0.00166f
C329 d4 comp_p_6/vinn 0.06841f
C330 comp_p_2/vinn comp_p_6/vbias_p 0.12413f
C331 d3 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C332 comp_p_6/vinn comp_p_6/latch_left 0.00473f
C333 comp_p_6/vbias_p comp_p_2/out_left 0.68901f
C334 d1 comp_p_3/latch_right 0
C335 d6 comp_p_3/latch_right 0.00265f
C336 d4 comp_p_4/vinn -0
C337 d5 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.00186f
C338 vbias_generation_0/XR_bias_3/R2 vdd 0.00793f
C339 d2 comp_p_1/out_left 0
C340 comp_p_6/tail vin 0
C341 d5 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0
C342 comp_p_1/latch_left comp_p_0/latch_right 0.02598f
C343 comp_p_1/latch_left d1 0.09502f
C344 comp_p_1/latch_left d6 0
C345 d0 tmux_7therm_to_3bin_0/R1/R1 0.00538f
C346 comp_p_2/latch_right comp_p_2/vinn 0
C347 comp_p_6/vbias_p comp_p_0/vinn 0.12305f
C348 comp_p_6/vbias_p comp_p_6/out_left -0.05299f
C349 comp_p_2/vinn comp_p_2/latch_left 0
C350 comp_p_6/vbias_p comp_p_1/out_left -0.065f
C351 d5 d1 0.26099f
C352 d5 d6 4.44886f
C353 vin comp_p_4/tail 0.01181f
C354 comp_p_1/vinn comp_p_0/latch_right 0.1958f
C355 d1 comp_p_1/vinn 0.26331f
C356 d6 comp_p_1/vinn 0
C357 d4 comp_p_6/latch_right 0.06065f
C358 d1 d0 1.12322f
C359 comp_p_2/latch_left comp_p_0/vinn 0
C360 d0 d6 0.09283f
C361 comp_p_5/vinn comp_p_5/latch_left 0.00674f
C362 vbias_generation_0/XR_bias_2/R2 vdd 0
C363 comp_p_6/vbias_p comp_p_5/out_left -0.0642f
C364 comp_p_6/vinn vbias_generation_0/XR_bias_4/R1 0.51064f
C365 comp_p_3/latch_left vdd 2.04611f
C366 comp_p_0/out_left vin 0.0787f
C367 d3 comp_p_3/vinn 0.0076f
C368 d2 comp_p_6/vbias_p 0.37534f
C369 d2 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C370 comp_p_0/latch_left comp_p_2/out_left 0.01472f
C371 d3 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C372 vbias_generation_0/bias_n comp_p_6/vinn 0.43753f
C373 comp_p_4/latch_right comp_p_6/vinn 0.00583f
C374 tmux_7therm_to_3bin_0/R1/R1 vdd 0.00399f
C375 vdd tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.00104f
C376 d4 comp_p_6/out_left 0.27385f
C377 d4 comp_p_1/out_left 0
C378 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vdd 0
C379 comp_p_4/latch_right comp_p_4/vinn 0.00144f
C380 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin vdd 0.00122f
C381 comp_p_0/latch_left comp_p_0/vinn 0.02494f
C382 comp_p_2/latch_right d2 0.00137f
C383 tmux_7therm_to_3bin_0/buffer_2/out d2 0
C384 d6 comp_p_5/latch_right 0
C385 comp_p_5/vinn comp_p_4/out_left 0.01843f
C386 comp_p_2/latch_right comp_p_6/vbias_p 0.40389f
C387 d1 vdd 1.15842f
C388 comp_p_0/latch_right vdd 0.00588f
C389 vin comp_p_0/tail 0.01181f
C390 d6 vdd 5.14819f
C391 comp_p_6/vbias_p comp_p_2/latch_left 0.37827f
C392 d4 comp_p_5/out_left 0.61081f
C393 d3 tmux_7therm_to_3bin_0/buffer_0/out 0
C394 d3 comp_p_1/latch_right 0.00104f
C395 comp_p_6/vinn vdd 0.76474f
C396 comp_p_1/vinn comp_p_2/out_left 0.00265f
C397 comp_p_5/vinn comp_p_3/vinn 0.0226f
C398 tmux_7therm_to_3bin_0/tmux_2to1_3/A vss 0.4939f
C399 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G vss 0.55051f
C400 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin vss 0.52606f
C401 dout2 vss 0.32356f
C402 tmux_7therm_to_3bin_0/buffer_8/inv_1/vin vss 0.52606f
C403 dout1 vss 0.32356f
C404 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vss 0.52606f
C405 dout0 vss 0.32356f
C406 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin vss 0.52765f
C407 tmux_7therm_to_3bin_0/buffer_6/out vss 0.67609f
C408 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin vss 0.52606f
C409 tmux_7therm_to_3bin_0/buffer_5/out vss 0.70857f
C410 vdd vss 0.37724p
C411 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vss 0.52606f
C412 tmux_7therm_to_3bin_0/buffer_4/out vss 0.70167f
C413 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin vss 0.52606f
C414 tmux_7therm_to_3bin_0/R1/R2 vss 0.22083f
C415 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin vss 0.52811f
C416 tmux_7therm_to_3bin_0/buffer_2/out vss 0.28552f
C417 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin vss 0.52606f
C418 tmux_7therm_to_3bin_0/buffer_1/out vss 0.30295f
C419 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin vss 0.52606f
C420 tmux_7therm_to_3bin_0/buffer_0/out vss 0.30577f
C421 tmux_7therm_to_3bin_0/R1/m1_n100_n100# vss 0.10692f
C422 tmux_7therm_to_3bin_0/buffer_8/in vss 1.28735f
C423 tmux_7therm_to_3bin_0/buffer_7/in vss 0.74661f
C424 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vss 0.55051f
C425 tmux_7therm_to_3bin_0/R1/R1 vss 3f
C426 tmux_7therm_to_3bin_0/tmux_2to1_3/B vss 0.41874f
C427 tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G vss 0.55051f
C428 tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G vss 0.55051f
C429 vin vss 21.46772f
C430 comp_p_6/tail vss 1.09633f
C431 comp_p_6/vbias_p vss 15.30121f
C432 d6 vss 4.91925f
C433 comp_p_6/latch_right vss 3.49411f
C434 comp_p_6/out_left vss 2.08951f
C435 comp_p_6/latch_left vss 3.68918f
C436 comp_p_5/tail vss 1.09613f
C437 d5 vss 3.00569f
C438 comp_p_5/latch_right vss 3.49805f
C439 comp_p_5/out_left vss 2.08667f
C440 comp_p_5/latch_left vss 3.68855f
C441 comp_p_4/tail vss 1.56897f
C442 d4 vss 9.43973f
C443 comp_p_4/latch_right vss 5.50989f
C444 comp_p_4/out_left vss 4.34925f
C445 comp_p_4/latch_left vss 6.03696f
C446 comp_p_3/tail vss 1.09611f
C447 d3 vss 2.71104f
C448 comp_p_3/latch_right vss 3.5009f
C449 comp_p_3/out_left vss 2.06137f
C450 comp_p_3/latch_left vss 3.68751f
C451 comp_p_2/tail vss 1.56898f
C452 d2 vss 7.1799f
C453 comp_p_2/latch_right vss 5.49653f
C454 comp_p_2/out_left vss 4.34035f
C455 comp_p_2/latch_left vss 6.03407f
C456 comp_p_0/tail vss 1.56897f
C457 d1 vss 7.38418f
C458 comp_p_0/latch_right vss 5.50255f
C459 comp_p_0/out_left vss 4.40824f
C460 comp_p_0/latch_left vss 6.03535f
C461 comp_p_1/tail vss 1.09611f
C462 d0 vss 2.80029f
C463 comp_p_1/latch_right vss 3.49227f
C464 comp_p_1/out_left vss 2.0627f
C465 comp_p_1/latch_left vss 3.68751f
C466 comp_p_0/vinn vss 5.97591f
C467 comp_p_2/vinn vss 4.36523f
C468 comp_p_3/vinn vss 7.39187f
C469 comp_p_4/vinn vss 4.39841f
C470 comp_p_5/vinn vss 7.08701f
C471 comp_p_6/vinn vss 8.48697f
C472 comp_p_1/vinn vss 8.08405f
C473 vref vss 4.63995f
C474 vbias_generation_0/bias_n vss 2.57801f
C475 vbias_generation_0/XR_bias_4/R1 vss 1.57005f
C476 vbias_generation_0/XR_bias_3/R2 vss 1.81091f
C477 vbias_generation_0/XR_bias_2/R2 vss 1.47453f
.ends

.subckt tt_um_tinyflash_extracted clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND
XflashADC_3bit_0 uo_out[0] uo_out[1] uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out
+ flashADC_3bit_0/vbias_generation_0/bias_n flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin flashADC_3bit_0/comp_p_3/latch_left
+ flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in
+ flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in
+ flashADC_3bit_0/comp_p_5/latch_left flashADC_3bit_0/vbias_generation_0/XR_bias_2/R2
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/m1_n100_n100# flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin
+ flashADC_3bit_0/comp_p_6/latch_left flashADC_3bit_0/comp_p_1/out_left flashADC_3bit_0/comp_p_6/tail
+ flashADC_3bit_0/comp_p_0/latch_right flashADC_3bit_0/comp_p_1/latch_right flashADC_3bit_0/comp_p_2/latch_right
+ flashADC_3bit_0/comp_p_3/latch_right flashADC_3bit_0/comp_p_3/tail flashADC_3bit_0/comp_p_4/latch_right
+ flashADC_3bit_0/comp_p_5/latch_right flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out flashADC_3bit_0/comp_p_4/out_left
+ flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_6/latch_right flashADC_3bit_0/comp_p_0/tail
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 flashADC_3bit_0/comp_p_2/latch_left
+ flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G
+ uo_out[4] flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G
+ flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out
+ flashADC_3bit_0/comp_p_0/out_left flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G flashADC_3bit_0/comp_p_6/vinn
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out uo_out[5] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin
+ flashADC_3bit_0/comp_p_4/tail flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/comp_p_0/latch_left
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin
+ uo_out[7] flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B
+ flashADC_3bit_0/comp_p_1/tail flashADC_3bit_0/comp_p_0/vinn ua[0] flashADC_3bit_0/comp_p_6/out_left
+ flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A flashADC_3bit_0/comp_p_1/latch_left
+ VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out uio_out[0] uo_out[6] uo_out[3]
+ flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_2/vinn ua[1] flashADC_3bit_0/comp_p_5/out_left
+ flashADC_3bit_0/vbias_generation_0/XR_bias_3/R2 uio_out[1] VGND flashADC_3bit_0/comp_p_3/out_left
+ flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit
X0 flashADC_3bit_0/comp_p_0/tail ua[0].t7 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X1 VDPWR flashADC_3bit_0/comp_p_4/out_left.t0 flashADC_3bit_0/comp_p_4/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X2 flashADC_3bit_0/comp_p_6/tail ua[0].t25 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X3 flashADC_3bit_0/comp_p_4/tail ua[0].t16 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X4 flashADC_3bit_0/comp_p_2/tail ua[0].t9 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X5 flashADC_3bit_0/comp_p_5/tail ua[0].t22 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X6 VDPWR flashADC_3bit_0/comp_p_6/out_left.t0 flashADC_3bit_0/comp_p_6/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X7 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin uo_out[6].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X8 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin uo_out[5].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X9 VDPWR flashADC_3bit_0/comp_p_2/out_left.t0 flashADC_3bit_0/comp_p_2/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X10 flashADC_3bit_0/comp_p_2/tail ua[0].t8 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X11 VDPWR flashADC_3bit_0/comp_p_6/out_left.t2 uio_out[1] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X12 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin uio_out[0].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X13 flashADC_3bit_0/comp_p_1/tail ua[0].t0 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X14 flashADC_3bit_0/comp_p_3/tail ua[0].t15 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X15 flashADC_3bit_0/comp_p_4/tail ua[0].t17 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X16 flashADC_3bit_0/comp_p_5/tail ua[0].t23 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X17 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin uio_out[1].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X18 flashADC_3bit_0/comp_p_1/tail ua[0].t1 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X19 flashADC_3bit_0/comp_p_3/out_left flashADC_3bit_0/comp_p_3/latch_left.t3 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X20 flashADC_3bit_0/comp_p_6/tail ua[0].t27 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X21 flashADC_3bit_0/comp_p_0/latch_left.t1 flashADC_3bit_0/comp_p_0/latch_left.t0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X22 flashADC_3bit_0/comp_p_6/tail ua[0].t26 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X23 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin uo_out[4].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X24 VDPWR flashADC_3bit_0/comp_p_4/out_left.t2 uo_out[7] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X25 flashADC_3bit_0/comp_p_4/tail ua[0].t18 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X26 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X27 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin uo_out[7].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X28 flashADC_3bit_0/comp_p_0/latch_right flashADC_3bit_0/comp_p_0/latch_left.t2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X29 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin uio_out[1].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X30 flashADC_3bit_0/comp_p_0/out_left flashADC_3bit_0/comp_p_0/latch_left.t3 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X31 flashADC_3bit_0/comp_p_0/tail ua[0].t4 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X32 flashADC_3bit_0/comp_p_1/tail ua[0].t2 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X33 flashADC_3bit_0/comp_p_2/tail ua[0].t11 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X34 VDPWR flashADC_3bit_0/comp_p_3/out_left.t0 flashADC_3bit_0/comp_p_3/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X35 flashADC_3bit_0/comp_p_3/tail ua[0].t14 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X36 flashADC_3bit_0/comp_p_4/tail ua[0].t19 flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X37 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin uo_out[6].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X38 flashADC_3bit_0/comp_p_0/tail ua[0].t5 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X39 flashADC_3bit_0/comp_p_1/tail ua[0].t3 flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X40 VDPWR flashADC_3bit_0/comp_p_2/out_left.t2 uo_out[5] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X41 VDPWR flashADC_3bit_0/comp_p_3/out_left.t2 uo_out[6] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X42 flashADC_3bit_0/comp_p_3/latch_left.t1 flashADC_3bit_0/comp_p_3/latch_left.t0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X43 flashADC_3bit_0/comp_p_6/tail ua[0].t24 flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X44 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin uio_out[0].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X45 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin uo_out[5].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X46 flashADC_3bit_0/comp_p_5/tail ua[0].t20 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X47 flashADC_3bit_0/comp_p_3/tail ua[0].t13 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X48 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin uo_out[7].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X49 VDPWR flashADC_3bit_0/comp_p_1/out_left.t0 flashADC_3bit_0/comp_p_1/out_left.t1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X50 flashADC_3bit_0/comp_p_3/latch_right flashADC_3bit_0/comp_p_3/latch_left.t2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X51 flashADC_3bit_0/comp_p_3/tail ua[0].t12 flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X52 VDPWR flashADC_3bit_0/comp_p_1/out_left.t2 uo_out[3] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X53 flashADC_3bit_0/comp_p_5/tail ua[0].t21 flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X54 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin uo_out[4].t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X55 flashADC_3bit_0/comp_p_0/tail ua[0].t6 flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X56 flashADC_3bit_0/comp_p_2/tail ua[0].t10 flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X57 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3].t1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
R0 VGND.n143 VGND.n14 167213
R1 VGND.n980 VGND.n14 110069
R2 VGND.n980 VGND.n979 75006.2
R3 VGND.n907 VGND.n906 28828.4
R4 VGND.n473 VGND.n16 15045.2
R5 VGND.n148 VGND.n144 13450.7
R6 VGND.n141 VGND.n138 13450.7
R7 VGND.n160 VGND.n137 13450.7
R8 VGND.n877 VGND.n864 12770.2
R9 VGND.n871 VGND.n865 12770.2
R10 VGND.n862 VGND.n857 12770.2
R11 VGND.n854 VGND.n851 12770.2
R12 VGND.n848 VGND.n844 12770.2
R13 VGND.n887 VGND.n886 12770.2
R14 VGND.n841 VGND.n260 12770.2
R15 VGND.n899 VGND.n898 12770.2
R16 VGND.n258 VGND.n254 12770.2
R17 VGND.n979 VGND.n978 12066.7
R18 VGND.n978 VGND.n15 12039.7
R19 VGND.n908 VGND.n907 11644.9
R20 VGND.n474 VGND.n473 11496.8
R21 VGND.n923 VGND.n920 10655.8
R22 VGND.n475 VGND.n251 6402.87
R23 VGND.n984 VGND.n8 5440.68
R24 VGND.n45 VGND.n35 5440.68
R25 VGND.n959 VGND.n33 5440.68
R26 VGND.n628 VGND.n279 5440.68
R27 VGND.n512 VGND.n318 5440.68
R28 VGND.n619 VGND.n280 5440.68
R29 VGND.n522 VGND.n319 5440.68
R30 VGND.n220 VGND.n169 5255.26
R31 VGND.n81 VGND.n69 5255.26
R32 VGND.n91 VGND.n70 5255.26
R33 VGND.n576 VGND.n296 5255.26
R34 VGND.n504 VGND.n341 5255.26
R35 VGND.n615 VGND.n292 5255.26
R36 VGND.n483 VGND.n342 5255.26
R37 VGND.n225 VGND.n166 5116.21
R38 VGND.n166 VGND.n135 5116.21
R39 VGND.n226 VGND.n225 5116.21
R40 VGND.n226 VGND.n135 5116.21
R41 VGND.n981 VGND.n980 4754.9
R42 VGND.n194 VGND.n172 4536.79
R43 VGND.n215 VGND.n172 4536.79
R44 VGND.n206 VGND.n184 4536.79
R45 VGND.n207 VGND.n206 4536.79
R46 VGND.n119 VGND.n77 4536.79
R47 VGND.n85 VGND.n77 4536.79
R48 VGND.n949 VGND.n46 4536.79
R49 VGND.n951 VGND.n46 4536.79
R50 VGND.n55 VGND.n52 4536.79
R51 VGND.n948 VGND.n55 4536.79
R52 VGND.n87 VGND.n86 4536.79
R53 VGND.n117 VGND.n87 4536.79
R54 VGND.n609 VGND.n303 4536.79
R55 VGND.n580 VGND.n303 4536.79
R56 VGND.n838 VGND.n265 4536.79
R57 VGND.n838 VGND.n266 4536.79
R58 VGND.n534 VGND.n348 4536.79
R59 VGND.n477 VGND.n348 4536.79
R60 VGND.n549 VGND.n329 4536.79
R61 VGND.n330 VGND.n329 4536.79
R62 VGND.n276 VGND.n264 4536.79
R63 VGND.n593 VGND.n264 4536.79
R64 VGND.n582 VGND.n581 4536.79
R65 VGND.n607 VGND.n582 4536.79
R66 VGND.n334 VGND.n331 4536.79
R67 VGND.n547 VGND.n334 4536.79
R68 VGND.n479 VGND.n478 4536.79
R69 VGND.n532 VGND.n479 4536.79
R70 VGND.n976 VGND.n16 4301.43
R71 VGND.n220 VGND.n7 4131.21
R72 VGND.n197 VGND.n196 4131.21
R73 VGND.n200 VGND.n199 4131.21
R74 VGND.n213 VGND.n175 4131.21
R75 VGND.n209 VGND.n182 4131.21
R76 VGND.n69 VGND.n68 4131.21
R77 VGND.n123 VGND.n40 4131.21
R78 VGND.n957 VGND.n41 4131.21
R79 VGND.n125 VGND.n65 4131.21
R80 VGND.n952 VGND.n39 4131.21
R81 VGND.n70 VGND.n32 4131.21
R82 VGND.n104 VGND.n72 4131.21
R83 VGND.n54 VGND.n38 4131.21
R84 VGND.n103 VGND.n71 4131.21
R85 VGND.n107 VGND.n36 4131.21
R86 VGND.n568 VGND.n296 4131.21
R87 VGND.n613 VGND.n284 4131.21
R88 VGND.n634 VGND.n285 4131.21
R89 VGND.n567 VGND.n299 4131.21
R90 VGND.n629 VGND.n283 4131.21
R91 VGND.n507 VGND.n341 4131.21
R92 VGND.n538 VGND.n323 4131.21
R93 VGND.n555 VGND.n324 4131.21
R94 VGND.n344 VGND.n315 4131.21
R95 VGND.n557 VGND.n316 4131.21
R96 VGND.n615 VGND.n294 4131.21
R97 VGND.n586 VGND.n298 4131.21
R98 VGND.n592 VGND.n282 4131.21
R99 VGND.n297 VGND.n275 4131.21
R100 VGND.n636 VGND.n277 4131.21
R101 VGND.n488 VGND.n342 4131.21
R102 VGND.n540 VGND.n339 4131.21
R103 VGND.n333 VGND.n322 4131.21
R104 VGND.n490 VGND.n343 4131.21
R105 VGND.n521 VGND.n320 4131.21
R106 VGND.n410 VGND.n409 4116.13
R107 VGND.n984 VGND.n7 3945.79
R108 VGND.n196 VGND.n187 3945.79
R109 VGND.n199 VGND.n197 3945.79
R110 VGND.n213 VGND.n173 3945.79
R111 VGND.n209 VGND.n175 3945.79
R112 VGND.n68 VGND.n35 3945.79
R113 VGND.n123 VGND.n73 3945.79
R114 VGND.n957 VGND.n40 3945.79
R115 VGND.n125 VGND.n63 3945.79
R116 VGND.n65 VGND.n39 3945.79
R117 VGND.n959 VGND.n32 3945.79
R118 VGND.n93 VGND.n72 3945.79
R119 VGND.n104 VGND.n38 3945.79
R120 VGND.n88 VGND.n71 3945.79
R121 VGND.n103 VGND.n36 3945.79
R122 VGND.n568 VGND.n279 3945.79
R123 VGND.n613 VGND.n300 3945.79
R124 VGND.n634 VGND.n284 3945.79
R125 VGND.n306 VGND.n299 3945.79
R126 VGND.n567 VGND.n283 3945.79
R127 VGND.n507 VGND.n318 3945.79
R128 VGND.n538 VGND.n345 3945.79
R129 VGND.n555 VGND.n323 3945.79
R130 VGND.n503 VGND.n344 3945.79
R131 VGND.n557 VGND.n315 3945.79
R132 VGND.n294 VGND.n280 3945.79
R133 VGND.n600 VGND.n298 3945.79
R134 VGND.n586 VGND.n282 3945.79
R135 VGND.n583 VGND.n297 3945.79
R136 VGND.n636 VGND.n275 3945.79
R137 VGND.n488 VGND.n319 3945.79
R138 VGND.n540 VGND.n338 3945.79
R139 VGND.n339 VGND.n322 3945.79
R140 VGND.n480 VGND.n343 3945.79
R141 VGND.n490 VGND.n320 3945.79
R142 VGND.n842 VGND.n841 3876.26
R143 VGND.n848 VGND.n842 3876.26
R144 VGND.n878 VGND.n862 3876.26
R145 VGND.n878 VGND.n877 3876.26
R146 VGND.n868 VGND.n865 3876.26
R147 VGND.n872 VGND.n864 3876.26
R148 VGND.n872 VGND.n871 3876.26
R149 VGND.n871 VGND.n870 3876.26
R150 VGND.n877 VGND.n876 3876.26
R151 VGND.n876 VGND.n865 3876.26
R152 VGND.n882 VGND.n851 3876.26
R153 VGND.n882 VGND.n857 3876.26
R154 VGND.n863 VGND.n857 3876.26
R155 VGND.n864 VGND.n863 3876.26
R156 VGND.n887 VGND.n849 3876.26
R157 VGND.n854 VGND.n849 3876.26
R158 VGND.n855 VGND.n854 3876.26
R159 VGND.n862 VGND.n855 3876.26
R160 VGND.n850 VGND.n844 3876.26
R161 VGND.n886 VGND.n850 3876.26
R162 VGND.n886 VGND.n885 3876.26
R163 VGND.n885 VGND.n851 3876.26
R164 VGND.n888 VGND.n848 3876.26
R165 VGND.n888 VGND.n887 3876.26
R166 VGND.n898 VGND.n896 3876.26
R167 VGND.n896 VGND.n260 3876.26
R168 VGND.n893 VGND.n260 3876.26
R169 VGND.n893 VGND.n844 3876.26
R170 VGND.n900 VGND.n258 3876.26
R171 VGND.n900 VGND.n899 3876.26
R172 VGND.n899 VGND.n259 3876.26
R173 VGND.n841 VGND.n259 3876.26
R174 VGND.n904 VGND.n254 3876.26
R175 VGND.n897 VGND.n254 3876.26
R176 VGND.n898 VGND.n897 3876.26
R177 VGND.n258 VGND.n253 3876.26
R178 VGND.n907 VGND.n251 3303.94
R179 VGND.n194 VGND.n187 3227.32
R180 VGND.n200 VGND.n184 3227.32
R181 VGND.n215 VGND.n173 3227.32
R182 VGND.n207 VGND.n182 3227.32
R183 VGND.n119 VGND.n73 3227.32
R184 VGND.n949 VGND.n41 3227.32
R185 VGND.n85 VGND.n63 3227.32
R186 VGND.n952 VGND.n951 3227.32
R187 VGND.n93 VGND.n86 3227.32
R188 VGND.n948 VGND.n54 3227.32
R189 VGND.n117 VGND.n88 3227.32
R190 VGND.n107 VGND.n52 3227.32
R191 VGND.n609 VGND.n300 3227.32
R192 VGND.n285 VGND.n265 3227.32
R193 VGND.n580 VGND.n306 3227.32
R194 VGND.n629 VGND.n266 3227.32
R195 VGND.n534 VGND.n345 3227.32
R196 VGND.n549 VGND.n324 3227.32
R197 VGND.n503 VGND.n477 3227.32
R198 VGND.n330 VGND.n316 3227.32
R199 VGND.n600 VGND.n581 3227.32
R200 VGND.n593 VGND.n592 3227.32
R201 VGND.n607 VGND.n583 3227.32
R202 VGND.n277 VGND.n276 3227.32
R203 VGND.n478 VGND.n338 3227.32
R204 VGND.n547 VGND.n333 3227.32
R205 VGND.n532 VGND.n480 3227.32
R206 VGND.n521 VGND.n331 3227.32
R207 VGND.n977 VGND.n976 2670.7
R208 VGND.n475 VGND.n474 2649.46
R209 VGND.n977 VGND.n14 2623.51
R210 VGND.n458 VGND.n455 2306.06
R211 VGND.n471 VGND.n455 2306.06
R212 VGND.n458 VGND.n456 2306.06
R213 VGND.n471 VGND.n456 2306.06
R214 VGND.n922 VGND.n243 2306.06
R215 VGND.n930 VGND.n243 2306.06
R216 VGND.n922 VGND.n244 2306.06
R217 VGND.n930 VGND.n244 2306.06
R218 VGND.n462 VGND.n461 2306.06
R219 VGND.n461 VGND.n454 2306.06
R220 VGND.n463 VGND.n462 2306.06
R221 VGND.n463 VGND.n454 2306.06
R222 VGND.n918 VGND.n19 2306.06
R223 VGND.n918 VGND.n20 2306.06
R224 VGND.n974 VGND.n19 2306.06
R225 VGND.n974 VGND.n20 2306.06
R226 VGND.n916 VGND.n910 2306.06
R227 VGND.n916 VGND.n911 2306.06
R228 VGND.n910 VGND.n18 2306.06
R229 VGND.n911 VGND.n18 2306.06
R230 VGND.n440 VGND.n351 2306.06
R231 VGND.n451 VGND.n351 2306.06
R232 VGND.n440 VGND.n352 2306.06
R233 VGND.n451 VGND.n352 2306.06
R234 VGND.n427 VGND.n358 2306.06
R235 VGND.n437 VGND.n358 2306.06
R236 VGND.n427 VGND.n359 2306.06
R237 VGND.n437 VGND.n359 2306.06
R238 VGND.n414 VGND.n381 2306.06
R239 VGND.n412 VGND.n381 2306.06
R240 VGND.n424 VGND.n366 2306.06
R241 VGND.n424 VGND.n367 2306.06
R242 VGND.n393 VGND.n383 2306.06
R243 VGND.n408 VGND.n383 2306.06
R244 VGND.n393 VGND.n384 2306.06
R245 VGND.n408 VGND.n384 2306.06
R246 VGND.n389 VGND.n387 2306.06
R247 VGND.n396 VGND.n387 2306.06
R248 VGND.n390 VGND.n389 2306.06
R249 VGND.n396 VGND.n390 2306.06
R250 VGND.n442 VGND.n355 2306.06
R251 VGND.n355 VGND.n350 2306.06
R252 VGND.n443 VGND.n442 2306.06
R253 VGND.n443 VGND.n350 2306.06
R254 VGND.n429 VGND.n364 2306.06
R255 VGND.n364 VGND.n357 2306.06
R256 VGND.n430 VGND.n429 2306.06
R257 VGND.n430 VGND.n357 2306.06
R258 VGND.n697 VGND.n679 2306.06
R259 VGND.n688 VGND.n679 2306.06
R260 VGND.n697 VGND.n680 2306.06
R261 VGND.n688 VGND.n680 2306.06
R262 VGND.n707 VGND.n669 2306.06
R263 VGND.n699 VGND.n669 2306.06
R264 VGND.n707 VGND.n670 2306.06
R265 VGND.n699 VGND.n670 2306.06
R266 VGND.n808 VGND.n804 2306.06
R267 VGND.n808 VGND.n805 2306.06
R268 VGND.n818 VGND.n664 2306.06
R269 VGND.n665 VGND.n664 2306.06
R270 VGND.n770 VGND.n744 2306.06
R271 VGND.n785 VGND.n744 2306.06
R272 VGND.n770 VGND.n745 2306.06
R273 VGND.n785 VGND.n745 2306.06
R274 VGND.n754 VGND.n751 2306.06
R275 VGND.n767 VGND.n751 2306.06
R276 VGND.n754 VGND.n752 2306.06
R277 VGND.n767 VGND.n752 2306.06
R278 VGND.n686 VGND.n677 2306.06
R279 VGND.n690 VGND.n686 2306.06
R280 VGND.n687 VGND.n677 2306.06
R281 VGND.n690 VGND.n687 2306.06
R282 VGND.n675 VGND.n667 2306.06
R283 VGND.n701 VGND.n675 2306.06
R284 VGND.n676 VGND.n667 2306.06
R285 VGND.n701 VGND.n676 2306.06
R286 VGND.n810 VGND.n722 2306.06
R287 VGND.n810 VGND.n726 2306.06
R288 VGND.n816 VGND.n711 2306.06
R289 VGND.n711 VGND.n666 2306.06
R290 VGND.n782 VGND.n778 2306.06
R291 VGND.n782 VGND.n779 2306.06
R292 VGND.n801 VGND.n728 2306.06
R293 VGND.n801 VGND.n729 2306.06
R294 VGND.n772 VGND.n747 2306.06
R295 VGND.n776 VGND.n747 2306.06
R296 VGND.n772 VGND.n748 2306.06
R297 VGND.n776 VGND.n748 2306.06
R298 VGND.n759 VGND.n758 2306.06
R299 VGND.n758 VGND.n750 2306.06
R300 VGND.n760 VGND.n759 2306.06
R301 VGND.n760 VGND.n750 2306.06
R302 VGND.n924 VGND.n247 2306.06
R303 VGND.n928 VGND.n247 2306.06
R304 VGND.n924 VGND.n248 2306.06
R305 VGND.n928 VGND.n248 2306.06
R306 VGND.n983 VGND.n982 2187.9
R307 VGND.n689 VGND.n251 2168.06
R308 VGND.n539 VGND.n317 1455.1
R309 VGND.n556 VGND.n321 1455.1
R310 VGND.n614 VGND.n278 1455.1
R311 VGND.n635 VGND.n281 1455.1
R312 VGND.n124 VGND.n34 1455.1
R313 VGND.n958 VGND.n37 1455.1
R314 VGND.n978 VGND.n977 1401.31
R315 VGND.n377 VGND.n376 1390.59
R316 VGND.n376 VGND.n372 1390.59
R317 VGND.n378 VGND.n375 1390.59
R318 VGND.n378 VGND.n371 1390.59
R319 VGND.n661 VGND.n657 1390.59
R320 VGND.n661 VGND.n651 1390.59
R321 VGND.n658 VGND.n656 1390.59
R322 VGND.n658 VGND.n650 1390.59
R323 VGND.n714 VGND.n710 1390.59
R324 VGND.n714 VGND.n713 1390.59
R325 VGND.n724 VGND.n723 1390.59
R326 VGND.n725 VGND.n724 1390.59
R327 VGND.n738 VGND.n737 1390.59
R328 VGND.n737 VGND.n733 1390.59
R329 VGND.n739 VGND.n736 1390.59
R330 VGND.n739 VGND.n732 1390.59
R331 VGND.n539 VGND.n340 1389.8
R332 VGND.n556 VGND.n317 1389.8
R333 VGND.n614 VGND.n295 1389.8
R334 VGND.n635 VGND.n278 1389.8
R335 VGND.n124 VGND.n66 1389.8
R336 VGND.n958 VGND.n34 1389.8
R337 VGND.n151 VGND.n148 1367.41
R338 VGND.n156 VGND.n138 1367.41
R339 VGND.n156 VGND.n144 1367.41
R340 VGND.n149 VGND.n144 1367.41
R341 VGND.n140 VGND.n137 1367.41
R342 VGND.n141 VGND.n140 1367.41
R343 VGND.n142 VGND.n141 1367.41
R344 VGND.n148 VGND.n142 1367.41
R345 VGND.n161 VGND.n160 1367.41
R346 VGND.n160 VGND.n159 1367.41
R347 VGND.n159 VGND.n138 1367.41
R348 VGND.n163 VGND.n137 1367.41
R349 VGND.n866 VGND 1333.46
R350 VGND.n909 VGND.n908 1320.82
R351 VGND.n920 VGND.n909 1320.82
R352 VGND.n173 VGND.n169 1309.47
R353 VGND.n178 VGND.n175 1309.47
R354 VGND.n178 VGND.n7 1309.47
R355 VGND.n182 VGND.n8 1309.47
R356 VGND.n201 VGND.n200 1309.47
R357 VGND.n201 VGND.n182 1309.47
R358 VGND.n197 VGND.n186 1309.47
R359 VGND.n186 VGND.n175 1309.47
R360 VGND.n190 VGND.n187 1309.47
R361 VGND.n190 VGND.n173 1309.47
R362 VGND.n81 VGND.n63 1309.47
R363 VGND.n67 VGND.n65 1309.47
R364 VGND.n68 VGND.n67 1309.47
R365 VGND.n952 VGND.n45 1309.47
R366 VGND.n953 VGND.n41 1309.47
R367 VGND.n953 VGND.n952 1309.47
R368 VGND.n64 VGND.n40 1309.47
R369 VGND.n65 VGND.n64 1309.47
R370 VGND.n74 VGND.n73 1309.47
R371 VGND.n74 VGND.n63 1309.47
R372 VGND.n102 VGND.n32 1309.47
R373 VGND.n103 VGND.n102 1309.47
R374 VGND.n91 VGND.n88 1309.47
R375 VGND.n107 VGND.n33 1309.47
R376 VGND.n94 VGND.n88 1309.47
R377 VGND.n94 VGND.n93 1309.47
R378 VGND.n105 VGND.n103 1309.47
R379 VGND.n105 VGND.n104 1309.47
R380 VGND.n108 VGND.n107 1309.47
R381 VGND.n108 VGND.n54 1309.47
R382 VGND.n576 VGND.n306 1309.47
R383 VGND.n569 VGND.n567 1309.47
R384 VGND.n569 VGND.n568 1309.47
R385 VGND.n629 VGND.n628 1309.47
R386 VGND.n630 VGND.n285 1309.47
R387 VGND.n630 VGND.n629 1309.47
R388 VGND.n566 VGND.n284 1309.47
R389 VGND.n567 VGND.n566 1309.47
R390 VGND.n305 VGND.n300 1309.47
R391 VGND.n306 VGND.n305 1309.47
R392 VGND.n504 VGND.n503 1309.47
R393 VGND.n508 VGND.n315 1309.47
R394 VGND.n508 VGND.n507 1309.47
R395 VGND.n512 VGND.n316 1309.47
R396 VGND.n551 VGND.n324 1309.47
R397 VGND.n551 VGND.n316 1309.47
R398 VGND.n325 VGND.n323 1309.47
R399 VGND.n325 VGND.n315 1309.47
R400 VGND.n502 VGND.n345 1309.47
R401 VGND.n503 VGND.n502 1309.47
R402 VGND.n294 VGND.n293 1309.47
R403 VGND.n293 VGND.n275 1309.47
R404 VGND.n583 VGND.n292 1309.47
R405 VGND.n619 VGND.n277 1309.47
R406 VGND.n601 VGND.n583 1309.47
R407 VGND.n601 VGND.n600 1309.47
R408 VGND.n587 VGND.n275 1309.47
R409 VGND.n587 VGND.n586 1309.47
R410 VGND.n591 VGND.n277 1309.47
R411 VGND.n592 VGND.n591 1309.47
R412 VGND.n491 VGND.n488 1309.47
R413 VGND.n491 VGND.n490 1309.47
R414 VGND.n483 VGND.n480 1309.47
R415 VGND.n522 VGND.n521 1309.47
R416 VGND.n485 VGND.n480 1309.47
R417 VGND.n485 VGND.n338 1309.47
R418 VGND.n490 VGND.n489 1309.47
R419 VGND.n489 VGND.n339 1309.47
R420 VGND.n521 VGND.n520 1309.47
R421 VGND.n520 VGND.n333 1309.47
R422 VGND.n906 VGND.n252 1157.81
R423 VGND.n895 VGND.n894 1157.81
R424 VGND.n894 VGND.n843 1157.81
R425 VGND.n884 VGND.n843 1157.81
R426 VGND.n884 VGND.n883 1157.81
R427 VGND.n883 VGND.n856 1157.81
R428 VGND.n856 VGND.n12 1157.81
R429 VGND.n533 VGND.n476 1136.73
R430 VGND.n533 VGND.n340 1136.73
R431 VGND.n548 VGND.n321 1136.73
R432 VGND.n548 VGND.n332 1136.73
R433 VGND.n608 VGND.n304 1136.73
R434 VGND.n608 VGND.n295 1136.73
R435 VGND.n281 VGND.n263 1136.73
R436 VGND.n839 VGND.n263 1136.73
R437 VGND.n118 VGND.n78 1136.73
R438 VGND.n118 VGND.n66 1136.73
R439 VGND.n950 VGND.n37 1136.73
R440 VGND.n950 VGND.n53 1136.73
R441 VGND.n981 VGND.n13 1136.71
R442 VGND.n152 VGND 1103.06
R443 VGND.n920 VGND.n919 1057.25
R444 VGND.n414 VGND.n375 915.471
R445 VGND.n419 VGND.n375 915.471
R446 VGND.n419 VGND.n377 915.471
R447 VGND.n377 VGND.n366 915.471
R448 VGND.n412 VGND.n371 915.471
R449 VGND.n421 VGND.n371 915.471
R450 VGND.n421 VGND.n372 915.471
R451 VGND.n372 VGND.n367 915.471
R452 VGND.n804 VGND.n656 915.471
R453 VGND.n822 VGND.n656 915.471
R454 VGND.n822 VGND.n657 915.471
R455 VGND.n818 VGND.n657 915.471
R456 VGND.n805 VGND.n650 915.471
R457 VGND.n824 VGND.n650 915.471
R458 VGND.n824 VGND.n651 915.471
R459 VGND.n665 VGND.n651 915.471
R460 VGND.n723 VGND.n722 915.471
R461 VGND.n723 VGND.n655 915.471
R462 VGND.n710 VGND.n655 915.471
R463 VGND.n816 VGND.n710 915.471
R464 VGND.n726 VGND.n725 915.471
R465 VGND.n725 VGND.n653 915.471
R466 VGND.n713 VGND.n653 915.471
R467 VGND.n713 VGND.n666 915.471
R468 VGND.n778 VGND.n736 915.471
R469 VGND.n794 VGND.n736 915.471
R470 VGND.n794 VGND.n738 915.471
R471 VGND.n738 VGND.n728 915.471
R472 VGND.n779 VGND.n732 915.471
R473 VGND.n796 VGND.n732 915.471
R474 VGND.n796 VGND.n733 915.471
R475 VGND.n733 VGND.n729 915.471
R476 VGND.n979 VGND.n13 880.169
R477 VGND.n154 VGND.n153 873.957
R478 VGND.n147 VGND.n145 873.957
R479 VGND.n139 VGND.n136 873.957
R480 VGND.n875 VGND.n874 829.741
R481 VGND.n867 VGND.n861 829.741
R482 VGND.n860 VGND.n858 829.741
R483 VGND.n880 VGND.n879 829.741
R484 VGND.n852 VGND.n847 829.741
R485 VGND.n891 VGND.n890 829.741
R486 VGND.n261 VGND.n257 829.741
R487 VGND.n889 VGND.n845 829.741
R488 VGND.n902 VGND.n901 829.741
R489 VGND.n840 VGND.n252 797.468
R490 VGND.n165 VGND.n164 768.378
R491 VGND.n332 VGND.n304 751.02
R492 VGND.n229 VGND.n228 705.365
R493 VGND.n158 VGND.n11 698.064
R494 VGND.n158 VGND.n157 698.064
R495 VGND.n157 VGND.n143 698.064
R496 VGND.n976 VGND.n975 665.898
R497 VGND.n903 VGND.n255 623.912
R498 VGND VGND.n255 619.196
R499 VGND.n228 VGND.n227 597.97
R500 VGND.n391 VGND.n249 560.645
R501 VGND.n395 VGND.n391 560.645
R502 VGND.n394 VGND.n382 560.645
R503 VGND.n409 VGND.n382 560.645
R504 VGND.n413 VGND.n410 560.645
R505 VGND.n413 VGND.n373 560.645
R506 VGND.n420 VGND.n373 560.645
R507 VGND.n420 VGND.n374 560.645
R508 VGND.n374 VGND.n365 560.645
R509 VGND.n425 VGND.n365 560.645
R510 VGND.n428 VGND.n356 560.645
R511 VGND.n438 VGND.n356 560.645
R512 VGND.n441 VGND.n349 560.645
R513 VGND.n452 VGND.n349 560.645
R514 VGND.n749 VGND.n250 560.645
R515 VGND.n768 VGND.n749 560.645
R516 VGND.n771 VGND.n746 560.645
R517 VGND.n784 VGND.n746 560.645
R518 VGND.n783 VGND.n777 560.645
R519 VGND.n777 VGND.n734 560.645
R520 VGND.n795 VGND.n734 560.645
R521 VGND.n795 VGND.n735 560.645
R522 VGND.n735 VGND.n727 560.645
R523 VGND.n802 VGND.n727 560.645
R524 VGND.n809 VGND.n803 560.645
R525 VGND.n803 VGND.n652 560.645
R526 VGND.n823 VGND.n652 560.645
R527 VGND.n823 VGND.n654 560.645
R528 VGND.n817 VGND.n654 560.645
R529 VGND.n817 VGND.n709 560.645
R530 VGND.n708 VGND.n668 560.645
R531 VGND.n700 VGND.n668 560.645
R532 VGND.n698 VGND.n678 560.645
R533 VGND.n689 VGND.n678 560.645
R534 VGND.n923 VGND.n245 560.645
R535 VGND.n929 VGND.n245 560.645
R536 VGND.n453 VGND.n246 560.645
R537 VGND.n472 VGND.n453 560.645
R538 VGND.n982 VGND.n981 500.092
R539 VGND.n198 VGND.n183 490.01
R540 VGND.n208 VGND.n183 490.01
R541 VGND.n208 VGND.n9 490.01
R542 VGND.n983 VGND.n9 490.01
R543 VGND.n223 VGND.n222 441.099
R544 VGND.n428 VGND.n425 376.13
R545 VGND.n784 VGND.n783 376.13
R546 VGND.n809 VGND.n802 376.13
R547 VGND.n709 VGND.n708 376.13
R548 VGND.n395 VGND.n394 369.033
R549 VGND.n441 VGND.n438 369.033
R550 VGND.n771 VGND.n768 369.033
R551 VGND.n700 VGND.n698 369.033
R552 VGND.n929 VGND.n246 369.033
R553 VGND.n895 VGND.n840 360.339
R554 VGND.n812 VGND.n811 343.154
R555 VGND.n165 VGND 334.683
R556 VGND.n195 VGND.n174 333.916
R557 VGND.n214 VGND.n174 333.916
R558 VGND.n214 VGND.n168 333.916
R559 VGND.n221 VGND.n168 333.916
R560 VGND.n224 VGND.n223 333.916
R561 VGND.n224 VGND.n10 333.916
R562 VGND.n982 VGND.n10 309.183
R563 VGND.n97 VGND.n89 294.776
R564 VGND.n482 VGND.n481 294.776
R565 VGND.n837 VGND.n267 294.776
R566 VGND.n585 VGND.n584 294.776
R567 VGND.n594 VGND.n590 294.776
R568 VGND.n610 VGND.n302 294.776
R569 VGND.n550 VGND.n328 294.776
R570 VGND.n535 VGND.n347 294.776
R571 VGND.n546 VGND.n545 294.776
R572 VGND.n205 VGND.n204 294.776
R573 VGND.n193 VGND.n171 294.776
R574 VGND.n50 VGND.n43 294.776
R575 VGND.n120 VGND.n76 294.776
R576 VGND.n947 VGND.n946 294.776
R577 VGND.n431 VGND.n430 292.5
R578 VGND.n430 VGND.n356 292.5
R579 VGND.n364 VGND 292.5
R580 VGND.n364 VGND.n356 292.5
R581 VGND.n444 VGND.n443 292.5
R582 VGND.n443 VGND.n349 292.5
R583 VGND.n355 VGND 292.5
R584 VGND.n355 VGND.n349 292.5
R585 VGND.n390 VGND 292.5
R586 VGND.n391 VGND.n390 292.5
R587 VGND.n387 VGND.n386 292.5
R588 VGND.n391 VGND.n387 292.5
R589 VGND VGND.n384 292.5
R590 VGND.n384 VGND.n382 292.5
R591 VGND.n385 VGND.n383 292.5
R592 VGND.n383 VGND.n382 292.5
R593 VGND VGND.n367 292.5
R594 VGND.n367 VGND.n365 292.5
R595 VGND VGND.n421 292.5
R596 VGND.n421 VGND.n420 292.5
R597 VGND.n412 VGND 292.5
R598 VGND.n413 VGND.n412 292.5
R599 VGND.n415 VGND.n414 292.5
R600 VGND.n414 VGND.n413 292.5
R601 VGND.n419 VGND.n418 292.5
R602 VGND.n420 VGND.n419 292.5
R603 VGND.n368 VGND.n366 292.5
R604 VGND.n366 VGND.n365 292.5
R605 VGND VGND.n359 292.5
R606 VGND.n359 VGND.n356 292.5
R607 VGND.n360 VGND.n358 292.5
R608 VGND.n358 VGND.n356 292.5
R609 VGND VGND.n352 292.5
R610 VGND.n352 VGND.n349 292.5
R611 VGND.n353 VGND.n351 292.5
R612 VGND.n351 VGND.n349 292.5
R613 VGND.n761 VGND.n760 292.5
R614 VGND.n760 VGND.n749 292.5
R615 VGND.n758 VGND 292.5
R616 VGND.n758 VGND.n749 292.5
R617 VGND.n774 VGND.n748 292.5
R618 VGND.n748 VGND.n746 292.5
R619 VGND VGND.n747 292.5
R620 VGND.n747 VGND.n746 292.5
R621 VGND.n799 VGND.n729 292.5
R622 VGND.n729 VGND.n727 292.5
R623 VGND.n797 VGND.n796 292.5
R624 VGND.n796 VGND.n795 292.5
R625 VGND.n780 VGND.n779 292.5
R626 VGND.n779 VGND.n777 292.5
R627 VGND VGND.n778 292.5
R628 VGND.n778 VGND.n777 292.5
R629 VGND.n794 VGND 292.5
R630 VGND.n795 VGND.n794 292.5
R631 VGND VGND.n728 292.5
R632 VGND.n728 VGND.n727 292.5
R633 VGND.n717 VGND.n666 292.5
R634 VGND.n817 VGND.n666 292.5
R635 VGND.n719 VGND.n653 292.5
R636 VGND.n823 VGND.n653 292.5
R637 VGND.n726 VGND.n721 292.5
R638 VGND.n803 VGND.n726 292.5
R639 VGND.n722 VGND 292.5
R640 VGND.n803 VGND.n722 292.5
R641 VGND VGND.n655 292.5
R642 VGND.n823 VGND.n655 292.5
R643 VGND.n816 VGND 292.5
R644 VGND.n817 VGND.n816 292.5
R645 VGND.n676 VGND.n674 292.5
R646 VGND.n676 VGND.n668 292.5
R647 VGND.n675 VGND 292.5
R648 VGND.n675 VGND.n668 292.5
R649 VGND.n687 VGND.n685 292.5
R650 VGND.n687 VGND.n678 292.5
R651 VGND.n686 VGND 292.5
R652 VGND.n686 VGND.n678 292.5
R653 VGND VGND.n752 292.5
R654 VGND.n752 VGND.n749 292.5
R655 VGND.n753 VGND.n751 292.5
R656 VGND.n751 VGND.n749 292.5
R657 VGND.n745 VGND 292.5
R658 VGND.n746 VGND.n745 292.5
R659 VGND.n744 VGND.n743 292.5
R660 VGND.n746 VGND.n744 292.5
R661 VGND.n665 VGND 292.5
R662 VGND.n817 VGND.n665 292.5
R663 VGND VGND.n824 292.5
R664 VGND.n824 VGND.n823 292.5
R665 VGND VGND.n805 292.5
R666 VGND.n805 VGND.n803 292.5
R667 VGND.n806 VGND.n804 292.5
R668 VGND.n804 VGND.n803 292.5
R669 VGND.n822 VGND.n821 292.5
R670 VGND.n823 VGND.n822 292.5
R671 VGND.n819 VGND.n818 292.5
R672 VGND.n818 VGND.n817 292.5
R673 VGND VGND.n670 292.5
R674 VGND.n670 VGND.n668 292.5
R675 VGND.n671 VGND.n669 292.5
R676 VGND.n669 VGND.n668 292.5
R677 VGND VGND.n680 292.5
R678 VGND.n680 VGND.n678 292.5
R679 VGND.n681 VGND.n679 292.5
R680 VGND.n679 VGND.n678 292.5
R681 VGND VGND.n18 292.5
R682 VGND.n975 VGND.n18 292.5
R683 VGND.n916 VGND.n915 292.5
R684 VGND.n919 VGND.n916 292.5
R685 VGND.n974 VGND 292.5
R686 VGND.n975 VGND.n974 292.5
R687 VGND.n918 VGND.n917 292.5
R688 VGND.n919 VGND.n918 292.5
R689 VGND.n464 VGND.n463 292.5
R690 VGND.n463 VGND.n453 292.5
R691 VGND.n461 VGND 292.5
R692 VGND.n461 VGND.n453 292.5
R693 VGND.n244 VGND 292.5
R694 VGND.n245 VGND.n244 292.5
R695 VGND.n243 VGND.n242 292.5
R696 VGND.n245 VGND.n243 292.5
R697 VGND VGND.n456 292.5
R698 VGND.n456 VGND.n453 292.5
R699 VGND.n457 VGND.n455 292.5
R700 VGND.n455 VGND.n453 292.5
R701 VGND.n926 VGND.n248 292.5
R702 VGND.n248 VGND.n245 292.5
R703 VGND VGND.n247 292.5
R704 VGND.n247 VGND.n245 292.5
R705 VGND VGND.n167 289.281
R706 VGND VGND.n134 285.604
R707 VGND.n621 VGND.n620 280.32
R708 VGND.n627 VGND.n626 280.32
R709 VGND.n514 VGND.n513 280.32
R710 VGND.n523 VGND.n519 280.32
R711 VGND.n985 VGND.n6 280.32
R712 VGND.n48 VGND.n47 280.32
R713 VGND.n960 VGND.n31 280.32
R714 VGND.n598 VGND.n597 268.425
R715 VGND.n596 VGND.n595 268.425
R716 VGND.n617 VGND.n616 268.425
R717 VGND.n575 VGND.n288 268.425
R718 VGND.n612 VGND.n286 268.425
R719 VGND.n633 VGND.n632 268.425
R720 VGND.n510 VGND.n506 268.425
R721 VGND.n537 VGND.n327 268.425
R722 VGND.n554 VGND.n553 268.425
R723 VGND.n494 VGND.n493 268.425
R724 VGND.n542 VGND.n541 268.425
R725 VGND.n544 VGND.n543 268.425
R726 VGND.n219 VGND.n5 268.425
R727 VGND.n189 VGND.n188 268.425
R728 VGND.n203 VGND.n185 268.425
R729 VGND.n80 VGND.n79 268.425
R730 VGND.n122 VGND.n42 268.425
R731 VGND.n956 VGND.n955 268.425
R732 VGND.n90 VGND.n30 268.425
R733 VGND.n101 VGND.n99 268.425
R734 VGND.n100 VGND.n56 268.425
R735 VGND.n616 VGND.n291 268.274
R736 VGND.n577 VGND.n575 268.274
R737 VGND.n506 VGND.n505 268.274
R738 VGND.n493 VGND.n484 268.274
R739 VGND.n219 VGND.n218 268.274
R740 VGND.n82 VGND.n80 268.274
R741 VGND.n92 VGND.n90 268.274
R742 VGND.n599 VGND.n598 256.377
R743 VGND.n597 VGND.n596 256.377
R744 VGND.n612 VGND.n611 256.377
R745 VGND.n633 VGND.n286 256.377
R746 VGND.n537 VGND.n536 256.377
R747 VGND.n554 VGND.n327 256.377
R748 VGND.n541 VGND.n337 256.377
R749 VGND.n543 VGND.n542 256.377
R750 VGND.n192 VGND.n189 256.377
R751 VGND.n188 VGND.n185 256.377
R752 VGND.n122 VGND.n121 256.377
R753 VGND.n956 VGND.n42 256.377
R754 VGND.n99 VGND.n98 256.377
R755 VGND.n101 VGND.n100 256.377
R756 VGND.n622 VGND.n621 256
R757 VGND.n626 VGND.n625 256
R758 VGND.n515 VGND.n514 256
R759 VGND.n519 VGND.n518 256
R760 VGND.n986 VGND.n985 256
R761 VGND.n47 VGND.n28 256
R762 VGND.n961 VGND.n960 256
R763 VGND.n902 VGND.n256 251.859
R764 VGND.n261 VGND.n256 251.859
R765 VGND.n853 VGND.n852 251.859
R766 VGND.n858 VGND.n853 251.859
R767 VGND.n874 VGND.n866 251.859
R768 VGND VGND.n861 251.859
R769 VGND VGND.n875 251.859
R770 VGND.n875 VGND 251.859
R771 VGND.n880 VGND.n859 251.859
R772 VGND.n867 VGND.n859 251.859
R773 VGND.n873 VGND.n867 251.859
R774 VGND.n874 VGND.n873 251.859
R775 VGND VGND.n860 251.859
R776 VGND.n879 VGND 251.859
R777 VGND.n879 VGND 251.859
R778 VGND VGND.n861 251.859
R779 VGND.n881 VGND.n858 251.859
R780 VGND.n881 VGND.n880 251.859
R781 VGND.n890 VGND 251.859
R782 VGND VGND.n847 251.859
R783 VGND VGND.n847 251.859
R784 VGND.n860 VGND 251.859
R785 VGND.n892 VGND.n845 251.859
R786 VGND.n892 VGND.n891 251.859
R787 VGND.n891 VGND.n846 251.859
R788 VGND.n852 VGND.n846 251.859
R789 VGND VGND.n257 251.859
R790 VGND.n889 VGND 251.859
R791 VGND VGND.n889 251.859
R792 VGND.n890 VGND 251.859
R793 VGND.n262 VGND.n261 251.859
R794 VGND.n845 VGND.n262 251.859
R795 VGND.n901 VGND 251.859
R796 VGND.n901 VGND 251.859
R797 VGND VGND.n257 251.859
R798 VGND.n903 VGND.n902 251.859
R799 VGND.n815 VGND.n814 249.667
R800 VGND.n599 VGND.n585 209.695
R801 VGND.n595 VGND.n594 209.695
R802 VGND.n611 VGND.n610 209.695
R803 VGND.n632 VGND.n267 209.695
R804 VGND.n536 VGND.n535 209.695
R805 VGND.n553 VGND.n550 209.695
R806 VGND.n481 VGND.n337 209.695
R807 VGND.n546 VGND.n544 209.695
R808 VGND.n193 VGND.n192 209.695
R809 VGND.n204 VGND.n203 209.695
R810 VGND.n121 VGND.n120 209.695
R811 VGND.n955 VGND.n43 209.695
R812 VGND.n98 VGND.n97 209.695
R813 VGND.n947 VGND.n56 209.695
R814 VGND.n909 VGND.n249 188.065
R815 VGND.n474 VGND.n452 188.065
R816 VGND.n908 VGND.n250 188.065
R817 VGND.n473 VGND.n472 188.065
R818 VGND.n982 VGND.n11 160.775
R819 VGND.n423 VGND.n368 150.417
R820 VGND.n819 VGND.n663 150.417
R821 VGND.n717 VGND.n712 150.417
R822 VGND.n800 VGND.n799 150.417
R823 VGND.n459 VGND.n457 149.835
R824 VGND.n470 VGND.n457 149.835
R825 VGND VGND.n459 149.835
R826 VGND.n921 VGND.n242 149.835
R827 VGND.n931 VGND.n242 149.835
R828 VGND.n921 VGND 149.835
R829 VGND.n460 VGND 149.835
R830 VGND.n464 VGND.n460 149.835
R831 VGND.n465 VGND.n464 149.835
R832 VGND.n439 VGND.n353 149.835
R833 VGND.n439 VGND 149.835
R834 VGND.n450 VGND.n353 149.835
R835 VGND.n426 VGND.n360 149.835
R836 VGND.n426 VGND 149.835
R837 VGND.n436 VGND.n360 149.835
R838 VGND.n415 VGND.n380 149.835
R839 VGND.n392 VGND.n385 149.835
R840 VGND.n392 VGND 149.835
R841 VGND.n407 VGND.n385 149.835
R842 VGND.n388 VGND.n386 149.835
R843 VGND.n388 VGND 149.835
R844 VGND.n397 VGND.n386 149.835
R845 VGND.n445 VGND.n444 149.835
R846 VGND.n444 VGND.n354 149.835
R847 VGND.n354 VGND 149.835
R848 VGND.n363 VGND 149.835
R849 VGND.n431 VGND.n363 149.835
R850 VGND.n432 VGND.n431 149.835
R851 VGND.n696 VGND.n681 149.835
R852 VGND.n696 VGND 149.835
R853 VGND.n682 VGND.n681 149.835
R854 VGND.n706 VGND.n671 149.835
R855 VGND.n706 VGND 149.835
R856 VGND.n672 VGND.n671 149.835
R857 VGND.n807 VGND.n806 149.835
R858 VGND.n769 VGND.n743 149.835
R859 VGND.n769 VGND 149.835
R860 VGND.n786 VGND.n743 149.835
R861 VGND.n755 VGND.n753 149.835
R862 VGND VGND.n755 149.835
R863 VGND.n766 VGND.n753 149.835
R864 VGND.n691 VGND.n685 149.835
R865 VGND.n685 VGND.n684 149.835
R866 VGND.n684 VGND 149.835
R867 VGND.n702 VGND.n674 149.835
R868 VGND.n674 VGND.n673 149.835
R869 VGND.n673 VGND 149.835
R870 VGND.n775 VGND.n774 149.835
R871 VGND.n774 VGND.n773 149.835
R872 VGND.n773 VGND 149.835
R873 VGND.n811 VGND.n721 149.835
R874 VGND.n781 VGND.n780 149.835
R875 VGND.n757 VGND 149.835
R876 VGND.n761 VGND.n757 149.835
R877 VGND.n762 VGND.n761 149.835
R878 VGND.n917 VGND.n21 149.835
R879 VGND VGND.n21 149.835
R880 VGND.n917 VGND.n22 149.835
R881 VGND.n915 VGND.n912 149.835
R882 VGND VGND.n912 149.835
R883 VGND.n915 VGND.n914 149.835
R884 VGND.n927 VGND.n926 149.835
R885 VGND.n926 VGND.n925 149.835
R886 VGND.n925 VGND 149.835
R887 VGND.n470 VGND.n469 149.459
R888 VGND.n932 VGND.n931 149.459
R889 VGND.n466 VGND.n465 149.459
R890 VGND.n450 VGND.n449 149.459
R891 VGND.n436 VGND.n435 149.459
R892 VGND.n407 VGND.n406 149.459
R893 VGND.n398 VGND.n397 149.459
R894 VGND.n446 VGND.n445 149.459
R895 VGND.n433 VGND.n432 149.459
R896 VGND.n695 VGND.n682 149.459
R897 VGND.n705 VGND.n672 149.459
R898 VGND.n787 VGND.n786 149.459
R899 VGND.n766 VGND.n765 149.459
R900 VGND.n692 VGND.n691 149.459
R901 VGND.n703 VGND.n702 149.459
R902 VGND.n775 VGND.n742 149.459
R903 VGND.n763 VGND.n762 149.459
R904 VGND.n973 VGND.n22 149.459
R905 VGND.n914 VGND.n913 149.459
R906 VGND.n927 VGND.n241 149.459
R907 VGND.n814 VGND.n813 132.8
R908 VGND.n800 VGND 132.129
R909 VGND.n423 VGND 132.127
R910 VGND VGND.n663 132.127
R911 VGND VGND.n380 130.802
R912 VGND.n807 VGND 130.802
R913 VGND.n781 VGND 130.802
R914 VGND VGND.n167 130.32
R915 VGND.n813 VGND.n812 120.001
R916 VGND VGND 118.966
R917 VGND.n228 VGND.n135 117.272
R918 VGND.n432 VGND.n357 117.001
R919 VGND.n438 VGND.n357 117.001
R920 VGND.n429 VGND.n363 117.001
R921 VGND.n429 VGND.n428 117.001
R922 VGND.n445 VGND.n350 117.001
R923 VGND.n452 VGND.n350 117.001
R924 VGND.n442 VGND.n354 117.001
R925 VGND.n442 VGND.n441 117.001
R926 VGND.n397 VGND.n396 117.001
R927 VGND.n396 VGND.n395 117.001
R928 VGND.n389 VGND.n388 117.001
R929 VGND.n389 VGND.n249 117.001
R930 VGND.n408 VGND.n407 117.001
R931 VGND.n409 VGND.n408 117.001
R932 VGND.n393 VGND.n392 117.001
R933 VGND.n394 VGND.n393 117.001
R934 VGND.n379 VGND.n378 117.001
R935 VGND.n378 VGND.n373 117.001
R936 VGND.n376 VGND.n369 117.001
R937 VGND.n376 VGND.n374 117.001
R938 VGND.n424 VGND.n423 117.001
R939 VGND.n425 VGND.n424 117.001
R940 VGND.n381 VGND.n380 117.001
R941 VGND.n410 VGND.n381 117.001
R942 VGND.n437 VGND.n436 117.001
R943 VGND.n438 VGND.n437 117.001
R944 VGND.n427 VGND.n426 117.001
R945 VGND.n428 VGND.n427 117.001
R946 VGND.n451 VGND.n450 117.001
R947 VGND.n452 VGND.n451 117.001
R948 VGND.n440 VGND.n439 117.001
R949 VGND.n441 VGND.n440 117.001
R950 VGND.n762 VGND.n750 117.001
R951 VGND.n768 VGND.n750 117.001
R952 VGND.n759 VGND.n757 117.001
R953 VGND.n759 VGND.n250 117.001
R954 VGND.n776 VGND.n775 117.001
R955 VGND.n784 VGND.n776 117.001
R956 VGND.n773 VGND.n772 117.001
R957 VGND.n772 VGND.n771 117.001
R958 VGND.n740 VGND.n739 117.001
R959 VGND.n739 VGND.n734 117.001
R960 VGND.n737 VGND.n730 117.001
R961 VGND.n737 VGND.n735 117.001
R962 VGND.n801 VGND.n800 117.001
R963 VGND.n802 VGND.n801 117.001
R964 VGND.n782 VGND.n781 117.001
R965 VGND.n783 VGND.n782 117.001
R966 VGND.n724 VGND.n716 117.001
R967 VGND.n724 VGND.n652 117.001
R968 VGND.n715 VGND.n714 117.001
R969 VGND.n714 VGND.n654 117.001
R970 VGND.n712 VGND.n711 117.001
R971 VGND.n711 VGND.n709 117.001
R972 VGND.n811 VGND.n810 117.001
R973 VGND.n810 VGND.n809 117.001
R974 VGND.n702 VGND.n701 117.001
R975 VGND.n701 VGND.n700 117.001
R976 VGND.n673 VGND.n667 117.001
R977 VGND.n708 VGND.n667 117.001
R978 VGND.n691 VGND.n690 117.001
R979 VGND.n690 VGND.n689 117.001
R980 VGND.n684 VGND.n677 117.001
R981 VGND.n698 VGND.n677 117.001
R982 VGND.n767 VGND.n766 117.001
R983 VGND.n768 VGND.n767 117.001
R984 VGND.n755 VGND.n754 117.001
R985 VGND.n754 VGND.n250 117.001
R986 VGND.n786 VGND.n785 117.001
R987 VGND.n785 VGND.n784 117.001
R988 VGND.n770 VGND.n769 117.001
R989 VGND.n771 VGND.n770 117.001
R990 VGND.n659 VGND.n658 117.001
R991 VGND.n658 VGND.n652 117.001
R992 VGND.n662 VGND.n661 117.001
R993 VGND.n661 VGND.n654 117.001
R994 VGND.n664 VGND.n663 117.001
R995 VGND.n709 VGND.n664 117.001
R996 VGND.n808 VGND.n807 117.001
R997 VGND.n809 VGND.n808 117.001
R998 VGND.n699 VGND.n672 117.001
R999 VGND.n700 VGND.n699 117.001
R1000 VGND.n707 VGND.n706 117.001
R1001 VGND.n708 VGND.n707 117.001
R1002 VGND.n688 VGND.n682 117.001
R1003 VGND.n689 VGND.n688 117.001
R1004 VGND.n697 VGND.n696 117.001
R1005 VGND.n698 VGND.n697 117.001
R1006 VGND.n486 VGND.n485 117.001
R1007 VGND.n485 VGND.n340 117.001
R1008 VGND.n523 VGND.n522 117.001
R1009 VGND.n522 VGND.n321 117.001
R1010 VGND.n520 VGND.n335 117.001
R1011 VGND.n520 VGND.n321 117.001
R1012 VGND.n492 VGND.n491 117.001
R1013 VGND.n491 VGND.n317 117.001
R1014 VGND.n489 VGND.n336 117.001
R1015 VGND.n489 VGND.n317 117.001
R1016 VGND.n545 VGND.n334 117.001
R1017 VGND.n334 VGND.n332 117.001
R1018 VGND.n482 VGND.n479 117.001
R1019 VGND.n479 VGND.n476 117.001
R1020 VGND.n484 VGND.n483 117.001
R1021 VGND.n483 VGND.n340 117.001
R1022 VGND.n602 VGND.n601 117.001
R1023 VGND.n601 VGND.n295 117.001
R1024 VGND.n620 VGND.n619 117.001
R1025 VGND.n619 VGND.n281 117.001
R1026 VGND.n591 VGND.n589 117.001
R1027 VGND.n591 VGND.n281 117.001
R1028 VGND.n293 VGND.n290 117.001
R1029 VGND.n293 VGND.n278 117.001
R1030 VGND.n588 VGND.n587 117.001
R1031 VGND.n587 VGND.n278 117.001
R1032 VGND.n590 VGND.n264 117.001
R1033 VGND.n839 VGND.n264 117.001
R1034 VGND.n584 VGND.n582 117.001
R1035 VGND.n582 VGND.n304 117.001
R1036 VGND.n292 VGND.n291 117.001
R1037 VGND.n295 VGND.n292 117.001
R1038 VGND.n502 VGND.n346 117.001
R1039 VGND.n502 VGND.n340 117.001
R1040 VGND.n552 VGND.n551 117.001
R1041 VGND.n551 VGND.n321 117.001
R1042 VGND.n329 VGND.n328 117.001
R1043 VGND.n332 VGND.n329 117.001
R1044 VGND.n326 VGND.n325 117.001
R1045 VGND.n325 VGND.n317 117.001
R1046 VGND.n509 VGND.n508 117.001
R1047 VGND.n508 VGND.n317 117.001
R1048 VGND.n513 VGND.n512 117.001
R1049 VGND.n512 VGND.n321 117.001
R1050 VGND.n505 VGND.n504 117.001
R1051 VGND.n504 VGND.n340 117.001
R1052 VGND.n348 VGND.n347 117.001
R1053 VGND.n476 VGND.n348 117.001
R1054 VGND.n305 VGND.n301 117.001
R1055 VGND.n305 VGND.n295 117.001
R1056 VGND.n631 VGND.n630 117.001
R1057 VGND.n630 VGND.n281 117.001
R1058 VGND.n838 VGND.n837 117.001
R1059 VGND.n839 VGND.n838 117.001
R1060 VGND.n566 VGND.n565 117.001
R1061 VGND.n566 VGND.n278 117.001
R1062 VGND.n570 VGND.n569 117.001
R1063 VGND.n569 VGND.n278 117.001
R1064 VGND.n628 VGND.n627 117.001
R1065 VGND.n628 VGND.n281 117.001
R1066 VGND.n577 VGND.n576 117.001
R1067 VGND.n576 VGND.n295 117.001
R1068 VGND.n303 VGND.n302 117.001
R1069 VGND.n304 VGND.n303 117.001
R1070 VGND.n95 VGND.n94 117.001
R1071 VGND.n94 VGND.n66 117.001
R1072 VGND.n33 VGND.n31 117.001
R1073 VGND.n37 VGND.n33 117.001
R1074 VGND.n109 VGND.n108 117.001
R1075 VGND.n108 VGND.n37 117.001
R1076 VGND.n102 VGND.n96 117.001
R1077 VGND.n102 VGND.n34 117.001
R1078 VGND.n106 VGND.n105 117.001
R1079 VGND.n105 VGND.n34 117.001
R1080 VGND.n946 VGND.n55 117.001
R1081 VGND.n55 VGND.n53 117.001
R1082 VGND.n89 VGND.n87 117.001
R1083 VGND.n87 VGND.n78 117.001
R1084 VGND.n92 VGND.n91 117.001
R1085 VGND.n91 VGND.n66 117.001
R1086 VGND.n75 VGND.n74 117.001
R1087 VGND.n74 VGND.n66 117.001
R1088 VGND.n954 VGND.n953 117.001
R1089 VGND.n953 VGND.n37 117.001
R1090 VGND.n50 VGND.n46 117.001
R1091 VGND.n53 VGND.n46 117.001
R1092 VGND.n64 VGND.n60 117.001
R1093 VGND.n64 VGND.n34 117.001
R1094 VGND.n67 VGND.n61 117.001
R1095 VGND.n67 VGND.n34 117.001
R1096 VGND.n48 VGND.n45 117.001
R1097 VGND.n45 VGND.n37 117.001
R1098 VGND.n82 VGND.n81 117.001
R1099 VGND.n81 VGND.n66 117.001
R1100 VGND.n77 VGND.n76 117.001
R1101 VGND.n78 VGND.n77 117.001
R1102 VGND.n164 VGND.n163 117.001
R1103 VGND.n146 VGND.n140 117.001
R1104 VGND.n158 VGND.n140 117.001
R1105 VGND VGND.n142 117.001
R1106 VGND.n157 VGND.n142 117.001
R1107 VGND.n152 VGND.n151 117.001
R1108 VGND.n149 VGND 117.001
R1109 VGND.n156 VGND.n155 117.001
R1110 VGND.n157 VGND.n156 117.001
R1111 VGND.n159 VGND 117.001
R1112 VGND.n159 VGND.n158 117.001
R1113 VGND.n161 VGND 117.001
R1114 VGND.n224 VGND.n135 117.001
R1115 VGND.n225 VGND 117.001
R1116 VGND.n225 VGND.n224 117.001
R1117 VGND.n191 VGND.n190 117.001
R1118 VGND.n190 VGND.n174 117.001
R1119 VGND.n186 VGND.n177 117.001
R1120 VGND.n186 VGND.n174 117.001
R1121 VGND.n179 VGND.n178 117.001
R1122 VGND.n178 VGND.n168 117.001
R1123 VGND.n218 VGND.n169 117.001
R1124 VGND.n169 VGND.n168 117.001
R1125 VGND.n172 VGND.n171 117.001
R1126 VGND.n174 VGND.n172 117.001
R1127 VGND.n202 VGND.n201 117.001
R1128 VGND.n201 VGND.n183 117.001
R1129 VGND.n206 VGND.n205 117.001
R1130 VGND.n206 VGND.n183 117.001
R1131 VGND.n8 VGND.n6 117.001
R1132 VGND.n9 VGND.n8 117.001
R1133 VGND.n914 VGND.n911 117.001
R1134 VGND.n911 VGND.n17 117.001
R1135 VGND.n912 VGND.n910 117.001
R1136 VGND.n910 VGND.n17 117.001
R1137 VGND.n22 VGND.n20 117.001
R1138 VGND.n20 VGND.n17 117.001
R1139 VGND.n21 VGND.n19 117.001
R1140 VGND.n19 VGND.n17 117.001
R1141 VGND.n465 VGND.n454 117.001
R1142 VGND.n472 VGND.n454 117.001
R1143 VGND.n462 VGND.n460 117.001
R1144 VGND.n462 VGND.n246 117.001
R1145 VGND.n931 VGND.n930 117.001
R1146 VGND.n930 VGND.n929 117.001
R1147 VGND.n922 VGND.n921 117.001
R1148 VGND.n923 VGND.n922 117.001
R1149 VGND.n471 VGND.n470 117.001
R1150 VGND.n472 VGND.n471 117.001
R1151 VGND.n459 VGND.n458 117.001
R1152 VGND.n458 VGND.n246 117.001
R1153 VGND.n928 VGND.n927 117.001
R1154 VGND.n929 VGND.n928 117.001
R1155 VGND.n925 VGND.n924 117.001
R1156 VGND.n924 VGND.n923 117.001
R1157 VGND VGND.n646 115.576
R1158 VGND.n151 VGND.n150 115.41
R1159 VGND.n162 VGND.n161 115.41
R1160 VGND.n163 VGND.n162 115.41
R1161 VGND.n150 VGND.n149 115.41
R1162 VGND.n476 VGND.n475 108.163
R1163 VGND.n840 VGND.n839 108.163
R1164 VGND.n78 VGND.n16 108.163
R1165 VGND.n222 VGND.n53 108.163
R1166 VGND.n167 VGND.n165 92.1893
R1167 VGND.n417 VGND.n369 90.3534
R1168 VGND.n422 VGND.n369 90.3534
R1169 VGND.n416 VGND.n379 90.3534
R1170 VGND.n411 VGND.n379 90.3534
R1171 VGND.n820 VGND.n662 90.3534
R1172 VGND.n662 VGND.n649 90.3534
R1173 VGND.n660 VGND.n659 90.3534
R1174 VGND.n659 VGND.n648 90.3534
R1175 VGND.n812 VGND.n716 90.3534
R1176 VGND.n720 VGND.n716 90.3534
R1177 VGND.n814 VGND.n715 90.3534
R1178 VGND.n718 VGND.n715 90.3534
R1179 VGND.n741 VGND.n740 90.3534
R1180 VGND.n740 VGND.n731 90.3534
R1181 VGND.n793 VGND.n730 90.3534
R1182 VGND.n798 VGND.n730 90.3534
R1183 VGND.n815 VGND.n712 89.9911
R1184 VGND.n154 VGND 88.8476
R1185 VGND VGND.n147 88.8476
R1186 VGND.n153 VGND 88.8476
R1187 VGND.n153 VGND.n152 88.8476
R1188 VGND VGND.n139 88.8476
R1189 VGND.n145 VGND 88.8476
R1190 VGND.n155 VGND.n145 88.8476
R1191 VGND.n155 VGND.n154 88.8476
R1192 VGND.n164 VGND.n136 88.8476
R1193 VGND.n146 VGND.n136 88.8476
R1194 VGND.n147 VGND.n146 88.8476
R1195 VGND.n139 VGND 88.8476
R1196 VGND.n597 VGND.n588 85.0829
R1197 VGND.n595 VGND.n589 85.0829
R1198 VGND.n602 VGND.n599 85.0829
R1199 VGND.n617 VGND.n290 85.0829
R1200 VGND.n290 VGND.n273 85.0829
R1201 VGND.n565 VGND.n286 85.0829
R1202 VGND.n572 VGND.n570 85.0829
R1203 VGND.n570 VGND.n288 85.0829
R1204 VGND.n611 VGND.n301 85.0829
R1205 VGND.n632 VGND.n631 85.0829
R1206 VGND.n327 VGND.n326 85.0829
R1207 VGND.n509 VGND.n313 85.0829
R1208 VGND.n510 VGND.n509 85.0829
R1209 VGND.n536 VGND.n346 85.0829
R1210 VGND.n553 VGND.n552 85.0829
R1211 VGND.n494 VGND.n492 85.0829
R1212 VGND.n527 VGND.n492 85.0829
R1213 VGND.n542 VGND.n336 85.0829
R1214 VGND.n544 VGND.n335 85.0829
R1215 VGND.n486 VGND.n337 85.0829
R1216 VGND.n188 VGND.n177 85.0829
R1217 VGND.n211 VGND.n179 85.0829
R1218 VGND.n179 VGND.n5 85.0829
R1219 VGND.n192 VGND.n191 85.0829
R1220 VGND.n203 VGND.n202 85.0829
R1221 VGND.n60 VGND.n42 85.0829
R1222 VGND.n127 VGND.n61 85.0829
R1223 VGND.n79 VGND.n61 85.0829
R1224 VGND.n121 VGND.n75 85.0829
R1225 VGND.n955 VGND.n954 85.0829
R1226 VGND.n96 VGND.n30 85.0829
R1227 VGND.n112 VGND.n96 85.0829
R1228 VGND.n106 VGND.n101 85.0829
R1229 VGND.n109 VGND.n56 85.0829
R1230 VGND.n98 VGND.n95 85.0829
R1231 VGND.n116 VGND.n89 84.9588
R1232 VGND.n531 VGND.n482 84.9588
R1233 VGND.n606 VGND.n584 84.9588
R1234 VGND.n579 VGND.n302 84.9588
R1235 VGND.n500 VGND.n347 84.9588
R1236 VGND.n216 VGND.n171 84.9588
R1237 VGND.n84 VGND.n76 84.9588
R1238 VGND.n837 VGND.n836 84.6953
R1239 VGND.n590 VGND.n269 84.6953
R1240 VGND.n328 VGND.n308 84.6953
R1241 VGND.n545 VGND.n309 84.6953
R1242 VGND.n205 VGND.n2 84.6953
R1243 VGND.n51 VGND.n50 84.6953
R1244 VGND.n946 VGND.n945 84.6953
R1245 VGND.n919 VGND.n17 83.7263
R1246 VGND.n975 VGND.n17 83.7263
R1247 VGND VGND.n815 77.2563
R1248 VGND.n222 VGND.n221 72.83
R1249 VGND.n603 VGND.n273 66.6518
R1250 VGND.n573 VGND.n572 66.6518
R1251 VGND.n498 VGND.n313 66.6518
R1252 VGND.n528 VGND.n527 66.6518
R1253 VGND.n212 VGND.n211 66.6518
R1254 VGND.n127 VGND.n126 66.6518
R1255 VGND.n113 VGND.n112 66.6518
R1256 VGND.n571 VGND.n287 64.7759
R1257 VGND.n637 VGND.n274 64.7759
R1258 VGND.n558 VGND.n314 64.7759
R1259 VGND.n526 VGND.n525 64.7759
R1260 VGND.n210 VGND.n181 64.7759
R1261 VGND.n128 VGND.n44 64.7759
R1262 VGND.n111 VGND.n110 64.7759
R1263 VGND.n572 VGND.n571 63.1207
R1264 VGND.n637 VGND.n273 63.1207
R1265 VGND.n558 VGND.n313 63.1207
R1266 VGND.n527 VGND.n526 63.1207
R1267 VGND.n211 VGND.n210 63.1207
R1268 VGND.n128 VGND.n127 63.1207
R1269 VGND.n112 VGND.n111 63.1207
R1270 VGND.n604 VGND.n603 61.2449
R1271 VGND.n574 VGND.n573 61.2449
R1272 VGND.n499 VGND.n498 61.2449
R1273 VGND.n529 VGND.n528 61.2449
R1274 VGND.n212 VGND.n170 61.2449
R1275 VGND.n126 VGND.n62 61.2449
R1276 VGND.n114 VGND.n113 61.2449
R1277 VGND.n416 VGND.n415 59.4829
R1278 VGND.n418 VGND.n416 59.4829
R1279 VGND.n418 VGND.n417 59.4829
R1280 VGND.n417 VGND.n368 59.4829
R1281 VGND.n806 VGND.n660 59.4829
R1282 VGND.n821 VGND.n660 59.4829
R1283 VGND.n821 VGND.n820 59.4829
R1284 VGND.n820 VGND.n819 59.4829
R1285 VGND.n721 VGND.n720 59.4829
R1286 VGND.n720 VGND.n719 59.4829
R1287 VGND.n719 VGND.n718 59.4829
R1288 VGND.n718 VGND.n717 59.4829
R1289 VGND.n780 VGND.n731 59.4829
R1290 VGND.n797 VGND.n731 59.4829
R1291 VGND.n798 VGND.n797 59.4829
R1292 VGND.n799 VGND.n798 59.4829
R1293 VGND.n589 VGND.n274 58.5793
R1294 VGND.n604 VGND.n602 58.5793
R1295 VGND.n574 VGND.n301 58.5793
R1296 VGND.n631 VGND.n287 58.5793
R1297 VGND.n499 VGND.n346 58.5793
R1298 VGND.n552 VGND.n314 58.5793
R1299 VGND.n525 VGND.n335 58.5793
R1300 VGND.n529 VGND.n486 58.5793
R1301 VGND.n191 VGND.n170 58.5793
R1302 VGND.n202 VGND.n181 58.5793
R1303 VGND.n75 VGND.n62 58.5793
R1304 VGND.n954 VGND.n44 58.5793
R1305 VGND.n110 VGND.n109 58.5793
R1306 VGND.n114 VGND.n95 58.5793
R1307 VGND.n588 VGND.n273 54.2123
R1308 VGND.n572 VGND.n565 54.2123
R1309 VGND.n326 VGND.n313 54.2123
R1310 VGND.n527 VGND.n336 54.2123
R1311 VGND.n211 VGND.n177 54.2123
R1312 VGND.n127 VGND.n60 54.2123
R1313 VGND.n112 VGND.n106 54.2123
R1314 VGND.n331 VGND.n309 41.7862
R1315 VGND.n548 VGND.n331 41.7862
R1316 VGND.n547 VGND.n546 41.7862
R1317 VGND.n548 VGND.n547 41.7862
R1318 VGND.n481 VGND.n478 41.7862
R1319 VGND.n533 VGND.n478 41.7862
R1320 VGND.n532 VGND.n531 41.7862
R1321 VGND.n533 VGND.n532 41.7862
R1322 VGND.n276 VGND.n269 41.7862
R1323 VGND.n276 VGND.n263 41.7862
R1324 VGND.n594 VGND.n593 41.7862
R1325 VGND.n593 VGND.n263 41.7862
R1326 VGND.n585 VGND.n581 41.7862
R1327 VGND.n608 VGND.n581 41.7862
R1328 VGND.n607 VGND.n606 41.7862
R1329 VGND.n608 VGND.n607 41.7862
R1330 VGND.n330 VGND.n308 41.7862
R1331 VGND.n548 VGND.n330 41.7862
R1332 VGND.n500 VGND.n477 41.7862
R1333 VGND.n533 VGND.n477 41.7862
R1334 VGND.n535 VGND.n534 41.7862
R1335 VGND.n534 VGND.n533 41.7862
R1336 VGND.n550 VGND.n549 41.7862
R1337 VGND.n549 VGND.n548 41.7862
R1338 VGND.n836 VGND.n266 41.7862
R1339 VGND.n266 VGND.n263 41.7862
R1340 VGND.n580 VGND.n579 41.7862
R1341 VGND.n608 VGND.n580 41.7862
R1342 VGND.n610 VGND.n609 41.7862
R1343 VGND.n609 VGND.n608 41.7862
R1344 VGND.n267 VGND.n265 41.7862
R1345 VGND.n265 VGND.n263 41.7862
R1346 VGND.n945 VGND.n52 41.7862
R1347 VGND.n950 VGND.n52 41.7862
R1348 VGND.n948 VGND.n947 41.7862
R1349 VGND.n950 VGND.n948 41.7862
R1350 VGND.n97 VGND.n86 41.7862
R1351 VGND.n118 VGND.n86 41.7862
R1352 VGND.n117 VGND.n116 41.7862
R1353 VGND.n118 VGND.n117 41.7862
R1354 VGND.n951 VGND.n51 41.7862
R1355 VGND.n951 VGND.n950 41.7862
R1356 VGND.n85 VGND.n84 41.7862
R1357 VGND.n118 VGND.n85 41.7862
R1358 VGND.n120 VGND.n119 41.7862
R1359 VGND.n119 VGND.n118 41.7862
R1360 VGND.n949 VGND.n43 41.7862
R1361 VGND.n950 VGND.n949 41.7862
R1362 VGND.n216 VGND.n215 41.7862
R1363 VGND.n215 VGND.n214 41.7862
R1364 VGND.n194 VGND.n193 41.7862
R1365 VGND.n195 VGND.n194 41.7862
R1366 VGND.n207 VGND.n2 41.7862
R1367 VGND.n208 VGND.n207 41.7862
R1368 VGND.n204 VGND.n184 41.7862
R1369 VGND.n198 VGND.n184 41.7862
R1370 VGND VGND.n411 40.4485
R1371 VGND.n422 VGND 40.4485
R1372 VGND VGND.n422 40.4485
R1373 VGND VGND.n648 40.4485
R1374 VGND VGND.n649 40.4485
R1375 VGND VGND.n649 40.4485
R1376 VGND VGND.n741 40.4485
R1377 VGND VGND.n793 40.4485
R1378 VGND.n793 VGND 40.4485
R1379 VGND.n411 VGND.n370 38.1445
R1380 VGND.n825 VGND.n648 38.1445
R1381 VGND.n792 VGND.n741 38.1445
R1382 VGND.n528 VGND.n343 34.4123
R1383 VGND.n539 VGND.n343 34.4123
R1384 VGND.n526 VGND.n320 34.4123
R1385 VGND.n556 VGND.n320 34.4123
R1386 VGND.n543 VGND.n322 34.4123
R1387 VGND.n556 VGND.n322 34.4123
R1388 VGND.n541 VGND.n540 34.4123
R1389 VGND.n540 VGND.n539 34.4123
R1390 VGND.n493 VGND.n342 34.4123
R1391 VGND.n539 VGND.n342 34.4123
R1392 VGND.n519 VGND.n319 34.4123
R1393 VGND.n556 VGND.n319 34.4123
R1394 VGND.n603 VGND.n297 34.4123
R1395 VGND.n614 VGND.n297 34.4123
R1396 VGND.n637 VGND.n636 34.4123
R1397 VGND.n636 VGND.n635 34.4123
R1398 VGND.n596 VGND.n282 34.4123
R1399 VGND.n635 VGND.n282 34.4123
R1400 VGND.n598 VGND.n298 34.4123
R1401 VGND.n614 VGND.n298 34.4123
R1402 VGND.n616 VGND.n615 34.4123
R1403 VGND.n615 VGND.n614 34.4123
R1404 VGND.n621 VGND.n280 34.4123
R1405 VGND.n635 VGND.n280 34.4123
R1406 VGND.n498 VGND.n344 34.4123
R1407 VGND.n539 VGND.n344 34.4123
R1408 VGND.n558 VGND.n557 34.4123
R1409 VGND.n557 VGND.n556 34.4123
R1410 VGND.n514 VGND.n318 34.4123
R1411 VGND.n556 VGND.n318 34.4123
R1412 VGND.n506 VGND.n341 34.4123
R1413 VGND.n539 VGND.n341 34.4123
R1414 VGND.n538 VGND.n537 34.4123
R1415 VGND.n539 VGND.n538 34.4123
R1416 VGND.n555 VGND.n554 34.4123
R1417 VGND.n556 VGND.n555 34.4123
R1418 VGND.n573 VGND.n299 34.4123
R1419 VGND.n614 VGND.n299 34.4123
R1420 VGND.n571 VGND.n283 34.4123
R1421 VGND.n635 VGND.n283 34.4123
R1422 VGND.n626 VGND.n279 34.4123
R1423 VGND.n635 VGND.n279 34.4123
R1424 VGND.n575 VGND.n296 34.4123
R1425 VGND.n614 VGND.n296 34.4123
R1426 VGND.n613 VGND.n612 34.4123
R1427 VGND.n614 VGND.n613 34.4123
R1428 VGND.n634 VGND.n633 34.4123
R1429 VGND.n635 VGND.n634 34.4123
R1430 VGND.n113 VGND.n71 34.4123
R1431 VGND.n124 VGND.n71 34.4123
R1432 VGND.n111 VGND.n36 34.4123
R1433 VGND.n958 VGND.n36 34.4123
R1434 VGND.n100 VGND.n38 34.4123
R1435 VGND.n958 VGND.n38 34.4123
R1436 VGND.n99 VGND.n72 34.4123
R1437 VGND.n124 VGND.n72 34.4123
R1438 VGND.n90 VGND.n70 34.4123
R1439 VGND.n124 VGND.n70 34.4123
R1440 VGND.n960 VGND.n959 34.4123
R1441 VGND.n959 VGND.n958 34.4123
R1442 VGND.n126 VGND.n125 34.4123
R1443 VGND.n125 VGND.n124 34.4123
R1444 VGND.n128 VGND.n39 34.4123
R1445 VGND.n958 VGND.n39 34.4123
R1446 VGND.n47 VGND.n35 34.4123
R1447 VGND.n958 VGND.n35 34.4123
R1448 VGND.n80 VGND.n69 34.4123
R1449 VGND.n124 VGND.n69 34.4123
R1450 VGND.n123 VGND.n122 34.4123
R1451 VGND.n124 VGND.n123 34.4123
R1452 VGND.n957 VGND.n956 34.4123
R1453 VGND.n958 VGND.n957 34.4123
R1454 VGND.n227 VGND.n226 34.4123
R1455 VGND.n226 VGND.n10 34.4123
R1456 VGND.n166 VGND.n134 34.4123
R1457 VGND.n223 VGND.n166 34.4123
R1458 VGND.n213 VGND.n212 34.4123
R1459 VGND.n214 VGND.n213 34.4123
R1460 VGND.n220 VGND.n219 34.4123
R1461 VGND.n221 VGND.n220 34.4123
R1462 VGND.n196 VGND.n189 34.4123
R1463 VGND.n196 VGND.n195 34.4123
R1464 VGND.n210 VGND.n209 34.4123
R1465 VGND.n209 VGND.n208 34.4123
R1466 VGND.n985 VGND.n984 34.4123
R1467 VGND.n984 VGND.n983 34.4123
R1468 VGND.n199 VGND.n185 34.4123
R1469 VGND.n199 VGND.n198 34.4123
R1470 VGND.n870 VGND.n866 32.5005
R1471 VGND.n876 VGND 32.5005
R1472 VGND.n876 VGND.n12 32.5005
R1473 VGND.n868 VGND 32.5005
R1474 VGND.n873 VGND.n872 32.5005
R1475 VGND.n872 VGND.n12 32.5005
R1476 VGND VGND.n878 32.5005
R1477 VGND.n878 VGND.n856 32.5005
R1478 VGND.n882 VGND.n881 32.5005
R1479 VGND.n883 VGND.n882 32.5005
R1480 VGND.n863 VGND.n859 32.5005
R1481 VGND.n863 VGND.n856 32.5005
R1482 VGND VGND.n855 32.5005
R1483 VGND.n883 VGND.n855 32.5005
R1484 VGND.n885 VGND.n853 32.5005
R1485 VGND.n885 VGND.n884 32.5005
R1486 VGND VGND.n888 32.5005
R1487 VGND.n888 VGND.n843 32.5005
R1488 VGND VGND.n849 32.5005
R1489 VGND.n884 VGND.n849 32.5005
R1490 VGND.n850 VGND.n846 32.5005
R1491 VGND.n850 VGND.n843 32.5005
R1492 VGND VGND.n842 32.5005
R1493 VGND.n894 VGND.n842 32.5005
R1494 VGND.n896 VGND.n262 32.5005
R1495 VGND.n896 VGND.n895 32.5005
R1496 VGND.n893 VGND.n892 32.5005
R1497 VGND.n894 VGND.n893 32.5005
R1498 VGND VGND.n259 32.5005
R1499 VGND.n895 VGND.n259 32.5005
R1500 VGND.n897 VGND.n256 32.5005
R1501 VGND.n897 VGND.n252 32.5005
R1502 VGND VGND.n253 32.5005
R1503 VGND VGND.n900 32.5005
R1504 VGND.n900 VGND.n252 32.5005
R1505 VGND.n904 VGND.n903 32.5005
R1506 VGND.n869 VGND.n868 32.3984
R1507 VGND.n870 VGND.n869 32.3984
R1508 VGND.n905 VGND.n904 32.3984
R1509 VGND.n905 VGND.n253 32.3984
R1510 VGND.n981 VGND.n12 21.0975
R1511 VGND.n618 VGND.n274 18.297
R1512 VGND.n605 VGND.n604 18.297
R1513 VGND.n578 VGND.n574 18.297
R1514 VGND.n287 VGND.n268 18.297
R1515 VGND.n501 VGND.n499 18.297
R1516 VGND.n511 VGND.n314 18.297
R1517 VGND.n525 VGND.n524 18.297
R1518 VGND.n530 VGND.n529 18.297
R1519 VGND.n217 VGND.n170 18.297
R1520 VGND.n181 VGND.n180 18.297
R1521 VGND.n83 VGND.n62 18.297
R1522 VGND.n49 VGND.n44 18.297
R1523 VGND.n110 VGND.n57 18.297
R1524 VGND.n115 VGND.n114 18.297
R1525 VGND.n116 VGND.n115 8.08353
R1526 VGND.n531 VGND.n530 8.08353
R1527 VGND.n606 VGND.n605 8.08353
R1528 VGND.n618 VGND.n269 8.08353
R1529 VGND.n579 VGND.n578 8.08353
R1530 VGND.n836 VGND.n268 8.08353
R1531 VGND.n501 VGND.n500 8.08353
R1532 VGND.n511 VGND.n308 8.08353
R1533 VGND.n524 VGND.n309 8.08353
R1534 VGND.n217 VGND.n216 8.08353
R1535 VGND.n180 VGND.n2 8.08353
R1536 VGND.n84 VGND.n83 8.08353
R1537 VGND.n51 VGND.n49 8.08353
R1538 VGND.n945 VGND.n57 8.08353
R1539 VGND.n969 VGND.n968 6.64112
R1540 VGND.n402 VGND.n362 5.57862
R1541 VGND.n828 VGND.n645 5.57706
R1542 VGND.n400 VGND 5.02361
R1543 VGND.n647 VGND 5.02361
R1544 VGND.n647 VGND 5.02361
R1545 VGND.n790 VGND 5.02361
R1546 VGND.n399 VGND 5.01717
R1547 VGND.n404 VGND 5.01717
R1548 VGND.n361 VGND 5.01717
R1549 VGND.n361 VGND 5.01717
R1550 VGND.n447 VGND 5.01717
R1551 VGND.n447 VGND 5.01717
R1552 VGND.n756 VGND 5.01717
R1553 VGND.n756 VGND 5.01717
R1554 VGND.n789 VGND 5.01717
R1555 VGND.n789 VGND 5.01717
R1556 VGND.n683 VGND 5.01717
R1557 VGND.n683 VGND 5.01717
R1558 VGND.n693 VGND 5.01717
R1559 VGND.n693 VGND 5.01717
R1560 VGND.n970 VGND 5.01717
R1561 VGND.n971 VGND 5.01717
R1562 VGND.n240 VGND 5.01717
R1563 VGND.n240 VGND 5.01717
R1564 VGND.n467 VGND 5.01717
R1565 VGND.n467 VGND 5.01717
R1566 VGND.n643 VGND 5.00093
R1567 VGND.n233 VGND 4.25376
R1568 VGND.n236 VGND 3.49683
R1569 VGND.n995 VGND 3.37909
R1570 VGND.n638 VGND.n272 3.27485
R1571 VGND.n559 VGND.n312 3.27485
R1572 VGND.n129 VGND.n26 3.27485
R1573 VGND.n58 VGND.n27 3.27485
R1574 VGND.n487 VGND.n310 3.27485
R1575 VGND.n564 VGND.n270 3.27485
R1576 VGND.n176 VGND.n3 3.27485
R1577 VGND.n620 VGND.n618 3.08756
R1578 VGND.n605 VGND.n291 3.08756
R1579 VGND.n578 VGND.n577 3.08756
R1580 VGND.n627 VGND.n268 3.08756
R1581 VGND.n505 VGND.n501 3.08756
R1582 VGND.n513 VGND.n511 3.08756
R1583 VGND.n524 VGND.n523 3.08756
R1584 VGND.n530 VGND.n484 3.08756
R1585 VGND.n218 VGND.n217 3.08756
R1586 VGND.n180 VGND.n6 3.08756
R1587 VGND.n83 VGND.n82 3.08756
R1588 VGND.n49 VGND.n48 3.08756
R1589 VGND.n57 VGND.n31 3.08756
R1590 VGND.n115 VGND.n92 3.08756
R1591 VGND.n307 VGND 3.06629
R1592 VGND.n496 VGND 3.06629
R1593 VGND.n964 VGND 3.06629
R1594 VGND.n813 VGND 3.01226
R1595 VGND.n640 VGND 2.51601
R1596 VGND.n935 VGND.n934 2.46929
R1597 VGND VGND.n370 2.3045
R1598 VGND.n825 VGND 2.3045
R1599 VGND VGND.n792 2.3045
R1600 VGND.n640 VGND 2.11902
R1601 VGND.n968 VGND.n24 1.98151
R1602 VGND.n399 VGND.n398 1.96988
R1603 VGND.n623 VGND 1.91991
R1604 VGND.n516 VGND 1.91991
R1605 VGND.n29 VGND 1.91991
R1606 VGND.n448 VGND.n446 1.8605
R1607 VGND.n406 VGND.n405 1.8605
R1608 VGND.n435 VGND.n434 1.8605
R1609 VGND.n449 VGND.n448 1.8605
R1610 VGND.n434 VGND.n433 1.8605
R1611 VGND.n788 VGND.n742 1.8605
R1612 VGND.n704 VGND.n703 1.8605
R1613 VGND.n694 VGND.n692 1.8605
R1614 VGND.n765 VGND.n764 1.8605
R1615 VGND.n788 VGND.n787 1.8605
R1616 VGND.n705 VGND.n704 1.8605
R1617 VGND.n695 VGND.n694 1.8605
R1618 VGND.n764 VGND.n763 1.8605
R1619 VGND.n913 VGND.n23 1.8605
R1620 VGND.n973 VGND.n972 1.8605
R1621 VGND.n933 VGND.n241 1.8605
R1622 VGND.n468 VGND.n466 1.8605
R1623 VGND.n933 VGND.n932 1.8605
R1624 VGND.n469 VGND.n468 1.8605
R1625 VGND.n829 VGND.n828 1.79344
R1626 VGND.n402 VGND.n235 1.68993
R1627 VGND.n130 VGND.n58 1.55665
R1628 VGND.n560 VGND.n310 1.55665
R1629 VGND.n639 VGND.n270 1.55665
R1630 VGND.n639 VGND.n638 1.55665
R1631 VGND.n560 VGND.n559 1.55665
R1632 VGND.n990 VGND.n3 1.55665
R1633 VGND.n130 VGND.n129 1.55665
R1634 VGND.n965 VGND.n27 1.43327
R1635 VGND.n495 VGND.n487 1.43327
R1636 VGND.n564 VGND.n563 1.43327
R1637 VGND.n563 VGND.n272 1.43327
R1638 VGND.n495 VGND.n312 1.43327
R1639 VGND.n176 VGND.n133 1.43327
R1640 VGND.n965 VGND.n26 1.43327
R1641 VGND.n229 VGND.n134 1.21955
R1642 VGND.n130 VGND 0.946224
R1643 VGND.n560 VGND 0.946224
R1644 VGND.n639 VGND 0.946224
R1645 VGND.n289 VGND 0.905763
R1646 VGND.n497 VGND 0.905763
R1647 VGND.n963 VGND 0.905763
R1648 VGND.n836 VGND.n835 0.846996
R1649 VGND.n835 VGND.n269 0.846996
R1650 VGND.n561 VGND.n308 0.846996
R1651 VGND.n561 VGND.n309 0.846996
R1652 VGND.n991 VGND.n2 0.846996
R1653 VGND.n944 VGND.n51 0.846996
R1654 VGND.n945 VGND.n944 0.846996
R1655 VGND VGND.n403 0.827844
R1656 VGND.n150 VGND.n143 0.796374
R1657 VGND.n162 VGND.n11 0.796374
R1658 VGND VGND 0.771099
R1659 VGND.n967 VGND.n25 0.760382
R1660 VGND.n401 VGND.n370 0.715885
R1661 VGND.n792 VGND.n791 0.715885
R1662 VGND.n826 VGND.n646 0.715885
R1663 VGND.n826 VGND.n825 0.715885
R1664 VGND.n988 VGND 0.695143
R1665 VGND.n571 VGND.n270 0.664786
R1666 VGND.n573 VGND.n564 0.664786
R1667 VGND.n638 VGND.n637 0.664786
R1668 VGND.n603 VGND.n272 0.664786
R1669 VGND.n559 VGND.n558 0.664786
R1670 VGND.n498 VGND.n312 0.664786
R1671 VGND.n526 VGND.n310 0.664786
R1672 VGND.n528 VGND.n487 0.664786
R1673 VGND.n210 VGND.n3 0.664786
R1674 VGND.n212 VGND.n176 0.664786
R1675 VGND.n231 VGND 0.664786
R1676 VGND.n129 VGND.n128 0.664786
R1677 VGND.n126 VGND.n26 0.664786
R1678 VGND.n111 VGND.n58 0.664786
R1679 VGND.n113 VGND.n27 0.664786
R1680 VGND.n4 VGND 0.644695
R1681 VGND.n644 VGND.n233 0.64299
R1682 VGND VGND 0.635531
R1683 VGND.n236 VGND.n234 0.629595
R1684 VGND.n227 VGND.n165 0.575781
R1685 VGND.n239 VGND.n24 0.568833
R1686 VGND.n238 VGND.n25 0.568833
R1687 VGND.n230 VGND.n229 0.517167
R1688 VGND VGND 0.457722
R1689 VGND.n59 VGND 0.447211
R1690 VGND.n311 VGND 0.447211
R1691 VGND.n271 VGND 0.447211
R1692 VGND.n563 VGND 0.439349
R1693 VGND.n495 VGND 0.439349
R1694 VGND.n965 VGND 0.439349
R1695 VGND VGND 0.406319
R1696 VGND.n791 VGND 0.405187
R1697 VGND.n827 VGND.n826 0.402844
R1698 VGND.n403 VGND.n401 0.401281
R1699 VGND.n562 VGND.n232 0.393625
R1700 VGND.n942 VGND.n941 0.393625
R1701 VGND.n469 VGND 0.376971
R1702 VGND.n932 VGND 0.376971
R1703 VGND.n466 VGND 0.376971
R1704 VGND.n449 VGND 0.376971
R1705 VGND.n435 VGND 0.376971
R1706 VGND.n406 VGND 0.376971
R1707 VGND.n398 VGND 0.376971
R1708 VGND.n446 VGND 0.376971
R1709 VGND.n433 VGND 0.376971
R1710 VGND VGND.n695 0.376971
R1711 VGND VGND.n705 0.376971
R1712 VGND.n787 VGND 0.376971
R1713 VGND.n765 VGND 0.376971
R1714 VGND.n692 VGND 0.376971
R1715 VGND.n703 VGND 0.376971
R1716 VGND VGND.n742 0.376971
R1717 VGND.n813 VGND.n646 0.376971
R1718 VGND.n763 VGND 0.376971
R1719 VGND.n622 VGND.n617 0.376971
R1720 VGND.n625 VGND.n288 0.376971
R1721 VGND.n515 VGND.n510 0.376971
R1722 VGND.n518 VGND.n494 0.376971
R1723 VGND.n986 VGND.n5 0.376971
R1724 VGND.n79 VGND.n28 0.376971
R1725 VGND VGND.n973 0.376971
R1726 VGND.n913 VGND 0.376971
R1727 VGND.n961 VGND.n30 0.376971
R1728 VGND VGND.n241 0.376971
R1729 VGND.n401 VGND.n400 0.376281
R1730 VGND.n791 VGND.n790 0.376281
R1731 VGND.n826 VGND.n647 0.376281
R1732 VGND.n238 VGND.n237 0.365484
R1733 VGND.n966 VGND.n965 0.346566
R1734 VGND.n990 VGND 0.342762
R1735 VGND.n59 VGND.n29 0.321553
R1736 VGND.n516 VGND.n311 0.321553
R1737 VGND.n623 VGND.n271 0.321553
R1738 VGND.n307 VGND.n289 0.321553
R1739 VGND.n497 VGND.n496 0.321553
R1740 VGND.n964 VGND.n963 0.321553
R1741 VGND.n989 VGND 0.318384
R1742 VGND.n642 VGND.n255 0.304262
R1743 VGND.n941 VGND.n940 0.285503
R1744 VGND.n643 VGND.n232 0.279901
R1745 VGND.n829 VGND.n235 0.250766
R1746 VGND.n935 VGND.n239 0.247336
R1747 VGND.n830 VGND 0.233324
R1748 VGND.n989 VGND.n988 0.228964
R1749 VGND.n642 VGND.n641 0.218382
R1750 VGND.n941 VGND.n0 0.209183
R1751 VGND.n972 VGND 0.208833
R1752 VGND VGND.n832 0.203416
R1753 VGND.n993 VGND.n1 0.203021
R1754 VGND.n936 VGND.n235 0.200936
R1755 VGND.n940 VGND.n232 0.196464
R1756 VGND.n641 VGND.n640 0.188289
R1757 VGND.n624 VGND.n289 0.186355
R1758 VGND.n517 VGND.n497 0.186355
R1759 VGND.n963 VGND.n962 0.186355
R1760 VGND.n834 VGND.n833 0.181262
R1761 VGND.n993 VGND.n992 0.181262
R1762 VGND.n130 VGND.n59 0.171553
R1763 VGND.n560 VGND.n311 0.171553
R1764 VGND.n639 VGND.n271 0.171553
R1765 VGND.n832 VGND.n642 0.169234
R1766 VGND.n943 VGND 0.166889
R1767 VGND.n434 VGND 0.166125
R1768 VGND.n704 VGND 0.166125
R1769 VGND.n405 VGND 0.164562
R1770 VGND.n448 VGND 0.164562
R1771 VGND.n788 VGND 0.164562
R1772 VGND.n694 VGND 0.164562
R1773 VGND.n468 VGND 0.164562
R1774 VGND.n624 VGND.n623 0.158395
R1775 VGND.n517 VGND.n516 0.158395
R1776 VGND.n962 VGND.n29 0.158395
R1777 VGND.n966 VGND.n23 0.14931
R1778 VGND.n563 VGND.n307 0.145237
R1779 VGND.n496 VGND.n495 0.145237
R1780 VGND.n965 VGND.n964 0.145237
R1781 VGND.n994 VGND.n993 0.144712
R1782 VGND.n972 VGND.n971 0.139389
R1783 VGND.n833 VGND.n1 0.137606
R1784 VGND.n624 VGND.n622 0.133357
R1785 VGND.n625 VGND.n624 0.133357
R1786 VGND.n517 VGND.n515 0.133357
R1787 VGND.n518 VGND.n517 0.133357
R1788 VGND.n987 VGND.n986 0.133357
R1789 VGND.n962 VGND.n28 0.133357
R1790 VGND.n962 VGND.n961 0.133357
R1791 VGND VGND.n4 0.126904
R1792 VGND.n937 VGND.n936 0.126796
R1793 VGND.n562 VGND 0.124938
R1794 VGND VGND.n943 0.123766
R1795 VGND.n641 VGND 0.111032
R1796 VGND.n969 VGND.n23 0.110619
R1797 VGND.n405 VGND.n404 0.109875
R1798 VGND.n448 VGND.n447 0.109875
R1799 VGND.n764 VGND.n756 0.109875
R1800 VGND.n789 VGND.n788 0.109875
R1801 VGND.n694 VGND.n693 0.109875
R1802 VGND.n468 VGND.n467 0.109875
R1803 VGND.n132 VGND 0.10256
R1804 VGND.n644 VGND 0.0991948
R1805 VGND.n434 VGND.n362 0.0934687
R1806 VGND.n967 VGND.n966 0.0907506
R1807 VGND.n704 VGND.n645 0.0903438
R1808 VGND.n934 VGND.n240 0.0860255
R1809 VGND.n234 VGND 0.0836655
R1810 VGND.n991 VGND.n990 0.0803611
R1811 VGND.n403 VGND.n402 0.0780862
R1812 VGND.n828 VGND.n827 0.0780862
R1813 VGND.n968 VGND.n967 0.0780862
R1814 VGND.n133 VGND 0.0759438
R1815 VGND VGND.n970 0.0699444
R1816 VGND.n971 VGND 0.0699444
R1817 VGND.n940 VGND.n939 0.0687
R1818 VGND VGND.n995 0.0686031
R1819 VGND.n987 VGND.n4 0.0677619
R1820 VGND.n835 VGND.n639 0.0651358
R1821 VGND.n561 VGND.n560 0.0651358
R1822 VGND VGND.n561 0.0651358
R1823 VGND.n944 VGND.n130 0.0651358
R1824 VGND.n944 VGND 0.0651358
R1825 VGND.n990 VGND.n989 0.0624048
R1826 VGND.n992 VGND 0.0620278
R1827 VGND.n988 VGND.n987 0.0576429
R1828 VGND.n834 VGND 0.0572671
R1829 VGND VGND.n399 0.0551875
R1830 VGND.n404 VGND 0.0551875
R1831 VGND.n361 VGND 0.0551875
R1832 VGND.n447 VGND 0.0551875
R1833 VGND.n756 VGND 0.0551875
R1834 VGND VGND.n789 0.0551875
R1835 VGND VGND.n683 0.0551875
R1836 VGND.n693 VGND 0.0551875
R1837 VGND VGND.n240 0.0551875
R1838 VGND.n467 VGND 0.0551875
R1839 VGND.n131 VGND 0.0524663
R1840 VGND.n869 VGND.n13 0.0523047
R1841 VGND.n906 VGND.n905 0.0523047
R1842 VGND.n936 VGND.n935 0.0501588
R1843 VGND.n938 VGND.n1 0.0478611
R1844 VGND.n400 VGND 0.0434688
R1845 VGND.n790 VGND 0.0434688
R1846 VGND VGND.n647 0.0434688
R1847 VGND.n131 VGND 0.0433241
R1848 VGND.n563 VGND.n562 0.042429
R1849 VGND.n132 VGND.n131 0.0417809
R1850 VGND.n133 VGND.n132 0.0416985
R1851 VGND VGND 0.0346797
R1852 VGND.n942 VGND.n231 0.0316884
R1853 VGND.n966 VGND 0.0297969
R1854 VGND.n943 VGND.n942 0.0294694
R1855 VGND.n970 VGND.n969 0.0292698
R1856 VGND.n934 VGND.n933 0.0233551
R1857 VGND.n683 VGND.n645 0.0200312
R1858 VGND.n992 VGND.n991 0.0188333
R1859 VGND.n362 VGND.n361 0.0169062
R1860 VGND.n832 VGND.n831 0.0134167
R1861 VGND.n230 VGND.n133 0.0120878
R1862 VGND.n239 VGND.n238 0.010792
R1863 VGND.n833 VGND 0.00952437
R1864 VGND.n835 VGND.n834 0.00836871
R1865 VGND VGND.n829 0.00513139
R1866 VGND.n25 VGND.n24 0.00492478
R1867 VGND.n827 VGND 0.00284375
R1868 VGND.n939 VGND.n233 0.00178858
R1869 VGND.n937 VGND.n234 0.00173884
R1870 VGND.n995 VGND.n994 0.00165108
R1871 VGND.n237 VGND.n236 0.00164397
R1872 VGND.n830 VGND.n644 0.00129115
R1873 VGND.n231 VGND.n230 0.000993097
R1874 VGND.n831 VGND.n830 0.00073924
R1875 VGND.n237 VGND.n0 0.000549738
R1876 VGND.n938 VGND.n937 0.000530793
R1877 VGND.n994 VGND.n0 0.000528422
R1878 VGND.n939 VGND.n938 0.00051895
R1879 VGND.n831 VGND.n643 0.000514212
R1880 VDPWR.n581 VDPWR.n577 5809.41
R1881 VDPWR.n624 VDPWR.n581 5809.41
R1882 VDPWR.n451 VDPWR.n340 5809.41
R1883 VDPWR.n340 VDPWR.n336 5809.41
R1884 VDPWR.n424 VDPWR.n360 5809.41
R1885 VDPWR.n424 VDPWR.n361 5809.41
R1886 VDPWR.n286 VDPWR.n138 5809.41
R1887 VDPWR.n286 VDPWR.n139 5809.41
R1888 VDPWR.n244 VDPWR.n145 5809.41
R1889 VDPWR.n163 VDPWR.n145 5809.41
R1890 VDPWR.n289 VDPWR.n288 5809.41
R1891 VDPWR.n288 VDPWR.n134 5809.41
R1892 VDPWR.n255 VDPWR.n146 5809.41
R1893 VDPWR.n255 VDPWR.n147 5809.41
R1894 VDPWR.n608 VDPWR.n605 5784.71
R1895 VDPWR.n609 VDPWR.n608 5784.71
R1896 VDPWR.n430 VDPWR.n429 5784.71
R1897 VDPWR.n429 VDPWR.n358 5784.71
R1898 VDPWR.n368 VDPWR.n365 5784.71
R1899 VDPWR.n419 VDPWR.n365 5784.71
R1900 VDPWR.n273 VDPWR.n268 5784.71
R1901 VDPWR.n269 VDPWR.n268 5784.71
R1902 VDPWR.n248 VDPWR.n157 5784.71
R1903 VDPWR.n157 VDPWR.n155 5784.71
R1904 VDPWR.n266 VDPWR.n257 5784.71
R1905 VDPWR.n266 VDPWR.n258 5784.71
R1906 VDPWR.n154 VDPWR.n151 5784.71
R1907 VDPWR.n250 VDPWR.n151 5784.71
R1908 VDPWR.n621 VDPWR.n584 4912.94
R1909 VDPWR.n621 VDPWR.n620 4912.94
R1910 VDPWR.n620 VDPWR.n585 4912.94
R1911 VDPWR.n585 VDPWR.n584 4912.94
R1912 VDPWR.n388 VDPWR.n384 4912.94
R1913 VDPWR.n400 VDPWR.n384 4912.94
R1914 VDPWR.n388 VDPWR.n385 4912.94
R1915 VDPWR.n400 VDPWR.n385 4912.94
R1916 VDPWR.n344 VDPWR.n343 4912.94
R1917 VDPWR.n448 VDPWR.n343 4912.94
R1918 VDPWR.n447 VDPWR.n344 4912.94
R1919 VDPWR.n448 VDPWR.n447 4912.94
R1920 VDPWR.n168 VDPWR.n165 4912.94
R1921 VDPWR.n241 VDPWR.n165 4912.94
R1922 VDPWR.n168 VDPWR.n166 4912.94
R1923 VDPWR.n241 VDPWR.n166 4912.94
R1924 VDPWR.n303 VDPWR.n120 4912.94
R1925 VDPWR.n282 VDPWR.n120 4912.94
R1926 VDPWR.n303 VDPWR.n121 4912.94
R1927 VDPWR.n282 VDPWR.n121 4912.94
R1928 VDPWR.n215 VDPWR.n193 4912.94
R1929 VDPWR.n215 VDPWR.n164 4912.94
R1930 VDPWR.n206 VDPWR.n193 4912.94
R1931 VDPWR.n206 VDPWR.n164 4912.94
R1932 VDPWR.n301 VDPWR.n123 4912.94
R1933 VDPWR.n280 VDPWR.n123 4912.94
R1934 VDPWR.n301 VDPWR.n124 4912.94
R1935 VDPWR.n280 VDPWR.n124 4912.94
R1936 VDPWR.n594 VDPWR.n593 4207.06
R1937 VDPWR.n576 VDPWR.n574 4207.06
R1938 VDPWR.n627 VDPWR.n574 4207.06
R1939 VDPWR.n617 VDPWR.n594 4207.06
R1940 VDPWR.n444 VDPWR.n348 4207.06
R1941 VDPWR.n348 VDPWR.n347 4207.06
R1942 VDPWR.n454 VDPWR.n333 4207.06
R1943 VDPWR.n335 VDPWR.n333 4207.06
R1944 VDPWR.n416 VDPWR.n372 4207.06
R1945 VDPWR.n372 VDPWR.n369 4207.06
R1946 VDPWR.n404 VDPWR.n377 4207.06
R1947 VDPWR.n383 VDPWR.n377 4207.06
R1948 VDPWR.n307 VDPWR.n111 4207.06
R1949 VDPWR.n309 VDPWR.n111 4207.06
R1950 VDPWR.n315 VDPWR.n107 4207.06
R1951 VDPWR.n107 VDPWR.n103 4207.06
R1952 VDPWR.n203 VDPWR.n202 4207.06
R1953 VDPWR.n202 VDPWR.n195 4207.06
R1954 VDPWR.n221 VDPWR.n220 4207.06
R1955 VDPWR.n222 VDPWR.n221 4207.06
R1956 VDPWR.n126 VDPWR.n116 4207.06
R1957 VDPWR.n126 VDPWR.n114 4207.06
R1958 VDPWR.n317 VDPWR.n101 4207.06
R1959 VDPWR.n104 VDPWR.n101 4207.06
R1960 VDPWR.n179 VDPWR.n171 4207.06
R1961 VDPWR.n232 VDPWR.n171 4207.06
R1962 VDPWR.n229 VDPWR.n173 4207.06
R1963 VDPWR.n230 VDPWR.n229 4207.06
R1964 VDPWR.n605 VDPWR.n597 4020
R1965 VDPWR.n609 VDPWR.n579 4020
R1966 VDPWR.n430 VDPWR.n338 4020
R1967 VDPWR.n358 VDPWR.n350 4020
R1968 VDPWR.n378 VDPWR.n368 4020
R1969 VDPWR.n419 VDPWR.n366 4020
R1970 VDPWR.n273 VDPWR.n272 4020
R1971 VDPWR.n270 VDPWR.n269 4020
R1972 VDPWR.n248 VDPWR.n158 4020
R1973 VDPWR.n211 VDPWR.n155 4020
R1974 VDPWR.n257 VDPWR.n133 4020
R1975 VDPWR.n260 VDPWR.n258 4020
R1976 VDPWR.n207 VDPWR.n154 4020
R1977 VDPWR.n250 VDPWR.n152 4020
R1978 VDPWR.n597 VDPWR.n577 3998.82
R1979 VDPWR.n624 VDPWR.n579 3998.82
R1980 VDPWR.n451 VDPWR.n338 3998.82
R1981 VDPWR.n350 VDPWR.n336 3998.82
R1982 VDPWR.n378 VDPWR.n360 3998.82
R1983 VDPWR.n366 VDPWR.n361 3998.82
R1984 VDPWR.n272 VDPWR.n138 3998.82
R1985 VDPWR.n270 VDPWR.n139 3998.82
R1986 VDPWR.n244 VDPWR.n158 3998.82
R1987 VDPWR.n211 VDPWR.n163 3998.82
R1988 VDPWR.n289 VDPWR.n133 3998.82
R1989 VDPWR.n260 VDPWR.n134 3998.82
R1990 VDPWR.n207 VDPWR.n146 3998.82
R1991 VDPWR.n152 VDPWR.n147 3998.82
R1992 VDPWR.n593 VDPWR.n592 3409.41
R1993 VDPWR.n592 VDPWR.n576 3409.41
R1994 VDPWR.n617 VDPWR.n573 3409.41
R1995 VDPWR.n627 VDPWR.n573 3409.41
R1996 VDPWR.n444 VDPWR.n332 3409.41
R1997 VDPWR.n454 VDPWR.n332 3409.41
R1998 VDPWR.n433 VDPWR.n347 3409.41
R1999 VDPWR.n433 VDPWR.n335 3409.41
R2000 VDPWR.n416 VDPWR.n373 3409.41
R2001 VDPWR.n404 VDPWR.n373 3409.41
R2002 VDPWR.n382 VDPWR.n369 3409.41
R2003 VDPWR.n383 VDPWR.n382 3409.41
R2004 VDPWR.n307 VDPWR.n106 3409.41
R2005 VDPWR.n315 VDPWR.n106 3409.41
R2006 VDPWR.n310 VDPWR.n309 3409.41
R2007 VDPWR.n310 VDPWR.n103 3409.41
R2008 VDPWR.n203 VDPWR.n187 3409.41
R2009 VDPWR.n220 VDPWR.n187 3409.41
R2010 VDPWR.n195 VDPWR.n186 3409.41
R2011 VDPWR.n222 VDPWR.n186 3409.41
R2012 VDPWR.n116 VDPWR.n100 3409.41
R2013 VDPWR.n317 VDPWR.n100 3409.41
R2014 VDPWR.n293 VDPWR.n114 3409.41
R2015 VDPWR.n293 VDPWR.n104 3409.41
R2016 VDPWR.n179 VDPWR.n178 3409.41
R2017 VDPWR.n178 VDPWR.n173 3409.41
R2018 VDPWR.n232 VDPWR.n231 3409.41
R2019 VDPWR.n231 VDPWR.n230 3409.41
R2020 VDPWR.n685 VDPWR.n670 1789.41
R2021 VDPWR.n692 VDPWR.n670 1789.41
R2022 VDPWR.n685 VDPWR.n671 1789.41
R2023 VDPWR.n692 VDPWR.n671 1789.41
R2024 VDPWR.n701 VDPWR.n663 1789.41
R2025 VDPWR.n682 VDPWR.n663 1789.41
R2026 VDPWR.n701 VDPWR.n664 1789.41
R2027 VDPWR.n682 VDPWR.n664 1789.41
R2028 VDPWR.n813 VDPWR.n806 1789.41
R2029 VDPWR.n806 VDPWR.n804 1789.41
R2030 VDPWR.n825 VDPWR.n658 1789.41
R2031 VDPWR.n827 VDPWR.n658 1789.41
R2032 VDPWR.n787 VDPWR.n768 1789.41
R2033 VDPWR.n787 VDPWR.n769 1789.41
R2034 VDPWR.n801 VDPWR.n727 1789.41
R2035 VDPWR.n801 VDPWR.n728 1789.41
R2036 VDPWR.n761 VDPWR.n733 1789.41
R2037 VDPWR.n790 VDPWR.n733 1789.41
R2038 VDPWR.n761 VDPWR.n734 1789.41
R2039 VDPWR.n790 VDPWR.n734 1789.41
R2040 VDPWR.n753 VDPWR.n745 1789.41
R2041 VDPWR.n745 VDPWR.n740 1789.41
R2042 VDPWR.n753 VDPWR.n746 1789.41
R2043 VDPWR.n746 VDPWR.n740 1789.41
R2044 VDPWR.n687 VDPWR.n673 1789.41
R2045 VDPWR.n690 VDPWR.n673 1789.41
R2046 VDPWR.n687 VDPWR.n674 1789.41
R2047 VDPWR.n690 VDPWR.n674 1789.41
R2048 VDPWR.n676 VDPWR.n661 1789.41
R2049 VDPWR.n681 VDPWR.n676 1789.41
R2050 VDPWR.n677 VDPWR.n661 1789.41
R2051 VDPWR.n681 VDPWR.n677 1789.41
R2052 VDPWR.n805 VDPWR.n724 1789.41
R2053 VDPWR.n815 VDPWR.n724 1789.41
R2054 VDPWR.n720 VDPWR.n704 1789.41
R2055 VDPWR.n720 VDPWR.n660 1789.41
R2056 VDPWR.n763 VDPWR.n736 1789.41
R2057 VDPWR.n766 VDPWR.n736 1789.41
R2058 VDPWR.n763 VDPWR.n737 1789.41
R2059 VDPWR.n766 VDPWR.n737 1789.41
R2060 VDPWR.n755 VDPWR.n741 1789.41
R2061 VDPWR.n758 VDPWR.n741 1789.41
R2062 VDPWR.n755 VDPWR.n742 1789.41
R2063 VDPWR.n758 VDPWR.n742 1789.41
R2064 VDPWR.n505 VDPWR.n479 1789.41
R2065 VDPWR.n479 VDPWR.n475 1789.41
R2066 VDPWR.n505 VDPWR.n480 1789.41
R2067 VDPWR.n480 VDPWR.n475 1789.41
R2068 VDPWR.n478 VDPWR.n472 1789.41
R2069 VDPWR.n507 VDPWR.n472 1789.41
R2070 VDPWR.n478 VDPWR.n473 1789.41
R2071 VDPWR.n507 VDPWR.n473 1789.41
R2072 VDPWR.n488 VDPWR.n483 1789.41
R2073 VDPWR.n497 VDPWR.n483 1789.41
R2074 VDPWR.n488 VDPWR.n484 1789.41
R2075 VDPWR.n497 VDPWR.n484 1789.41
R2076 VDPWR.n490 VDPWR.n486 1789.41
R2077 VDPWR.n495 VDPWR.n490 1789.41
R2078 VDPWR.n491 VDPWR.n486 1789.41
R2079 VDPWR.n495 VDPWR.n491 1789.41
R2080 VDPWR.n553 VDPWR.n527 1789.41
R2081 VDPWR.n527 VDPWR.n523 1789.41
R2082 VDPWR.n553 VDPWR.n528 1789.41
R2083 VDPWR.n528 VDPWR.n523 1789.41
R2084 VDPWR.n526 VDPWR.n520 1789.41
R2085 VDPWR.n555 VDPWR.n520 1789.41
R2086 VDPWR.n526 VDPWR.n521 1789.41
R2087 VDPWR.n555 VDPWR.n521 1789.41
R2088 VDPWR.n536 VDPWR.n531 1789.41
R2089 VDPWR.n545 VDPWR.n531 1789.41
R2090 VDPWR.n536 VDPWR.n532 1789.41
R2091 VDPWR.n545 VDPWR.n532 1789.41
R2092 VDPWR.n538 VDPWR.n534 1789.41
R2093 VDPWR.n543 VDPWR.n538 1789.41
R2094 VDPWR.n539 VDPWR.n534 1789.41
R2095 VDPWR.n543 VDPWR.n539 1789.41
R2096 VDPWR.n599 VDPWR.n597 1789.41
R2097 VDPWR.n599 VDPWR.n579 1789.41
R2098 VDPWR.n354 VDPWR.n338 1789.41
R2099 VDPWR.n354 VDPWR.n350 1789.41
R2100 VDPWR.n379 VDPWR.n378 1789.41
R2101 VDPWR.n379 VDPWR.n366 1789.41
R2102 VDPWR.n82 VDPWR.n5 1789.41
R2103 VDPWR.n85 VDPWR.n5 1789.41
R2104 VDPWR.n83 VDPWR.n82 1789.41
R2105 VDPWR.n76 VDPWR.n9 1789.41
R2106 VDPWR.n79 VDPWR.n9 1789.41
R2107 VDPWR.n76 VDPWR.n10 1789.41
R2108 VDPWR.n79 VDPWR.n10 1789.41
R2109 VDPWR.n56 VDPWR.n27 1789.41
R2110 VDPWR.n54 VDPWR.n27 1789.41
R2111 VDPWR.n73 VDPWR.n14 1789.41
R2112 VDPWR.n73 VDPWR.n15 1789.41
R2113 VDPWR.n48 VDPWR.n29 1789.41
R2114 VDPWR.n51 VDPWR.n29 1789.41
R2115 VDPWR.n48 VDPWR.n30 1789.41
R2116 VDPWR.n51 VDPWR.n30 1789.41
R2117 VDPWR.n45 VDPWR.n34 1789.41
R2118 VDPWR.n42 VDPWR.n35 1789.41
R2119 VDPWR.n45 VDPWR.n35 1789.41
R2120 VDPWR.n272 VDPWR.n271 1789.41
R2121 VDPWR.n271 VDPWR.n270 1789.41
R2122 VDPWR.n212 VDPWR.n158 1789.41
R2123 VDPWR.n212 VDPWR.n211 1789.41
R2124 VDPWR.n261 VDPWR.n133 1789.41
R2125 VDPWR.n261 VDPWR.n260 1789.41
R2126 VDPWR.n208 VDPWR.n207 1789.41
R2127 VDPWR.n208 VDPWR.n152 1789.41
R2128 VDPWR.n53 VDPWR.n52 1315.04
R2129 VDPWR.n706 VDPWR.n705 1231.76
R2130 VDPWR.n705 VDPWR.n657 1231.76
R2131 VDPWR.n808 VDPWR.n708 1231.76
R2132 VDPWR.n808 VDPWR.n807 1231.76
R2133 VDPWR.n777 VDPWR.n776 1231.76
R2134 VDPWR.n776 VDPWR.n775 1231.76
R2135 VDPWR.n782 VDPWR.n771 1231.76
R2136 VDPWR.n782 VDPWR.n772 1231.76
R2137 VDPWR.n716 VDPWR.n713 1231.76
R2138 VDPWR.n716 VDPWR.n715 1231.76
R2139 VDPWR.n817 VDPWR.n712 1231.76
R2140 VDPWR.n817 VDPWR.n816 1231.76
R2141 VDPWR.n25 VDPWR.n24 1231.76
R2142 VDPWR.n24 VDPWR.n20 1231.76
R2143 VDPWR.n58 VDPWR.n23 1231.76
R2144 VDPWR.n58 VDPWR.n19 1231.76
R2145 VDPWR.n592 VDPWR.n591 797.648
R2146 VDPWR.n591 VDPWR.n573 797.648
R2147 VDPWR.n434 VDPWR.n332 797.648
R2148 VDPWR.n434 VDPWR.n433 797.648
R2149 VDPWR.n381 VDPWR.n373 797.648
R2150 VDPWR.n382 VDPWR.n381 797.648
R2151 VDPWR.n311 VDPWR.n106 797.648
R2152 VDPWR.n311 VDPWR.n310 797.648
R2153 VDPWR.n210 VDPWR.n187 797.648
R2154 VDPWR.n210 VDPWR.n186 797.648
R2155 VDPWR.n294 VDPWR.n100 797.648
R2156 VDPWR.n294 VDPWR.n293 797.648
R2157 VDPWR.n178 VDPWR.n172 797.648
R2158 VDPWR.n231 VDPWR.n172 797.648
R2159 VDPWR.n813 VDPWR.n708 557.648
R2160 VDPWR.n823 VDPWR.n708 557.648
R2161 VDPWR.n823 VDPWR.n706 557.648
R2162 VDPWR.n825 VDPWR.n706 557.648
R2163 VDPWR.n807 VDPWR.n804 557.648
R2164 VDPWR.n807 VDPWR.n710 557.648
R2165 VDPWR.n710 VDPWR.n657 557.648
R2166 VDPWR.n827 VDPWR.n657 557.648
R2167 VDPWR.n771 VDPWR.n768 557.648
R2168 VDPWR.n779 VDPWR.n771 557.648
R2169 VDPWR.n779 VDPWR.n777 557.648
R2170 VDPWR.n777 VDPWR.n727 557.648
R2171 VDPWR.n772 VDPWR.n769 557.648
R2172 VDPWR.n773 VDPWR.n772 557.648
R2173 VDPWR.n775 VDPWR.n773 557.648
R2174 VDPWR.n775 VDPWR.n728 557.648
R2175 VDPWR.n805 VDPWR.n712 557.648
R2176 VDPWR.n821 VDPWR.n712 557.648
R2177 VDPWR.n821 VDPWR.n713 557.648
R2178 VDPWR.n713 VDPWR.n704 557.648
R2179 VDPWR.n816 VDPWR.n815 557.648
R2180 VDPWR.n816 VDPWR.n711 557.648
R2181 VDPWR.n715 VDPWR.n711 557.648
R2182 VDPWR.n715 VDPWR.n660 557.648
R2183 VDPWR.n56 VDPWR.n23 557.648
R2184 VDPWR.n68 VDPWR.n23 557.648
R2185 VDPWR.n68 VDPWR.n25 557.648
R2186 VDPWR.n25 VDPWR.n14 557.648
R2187 VDPWR.n54 VDPWR.n19 557.648
R2188 VDPWR.n70 VDPWR.n19 557.648
R2189 VDPWR.n70 VDPWR.n20 557.648
R2190 VDPWR.n20 VDPWR.n15 557.648
R2191 VDPWR.n602 VDPWR.n601 447.06
R2192 VDPWR.n352 VDPWR.n351 447.06
R2193 VDPWR.n423 VDPWR.n422 447.06
R2194 VDPWR.n245 VDPWR.n161 447.06
R2195 VDPWR.n285 VDPWR.n276 447.06
R2196 VDPWR.n259 VDPWR.n136 447.06
R2197 VDPWR.n254 VDPWR.n253 447.06
R2198 VDPWR.n604 VDPWR.n595 444.515
R2199 VDPWR.n357 VDPWR.n349 444.515
R2200 VDPWR.n420 VDPWR.n364 444.515
R2201 VDPWR.n247 VDPWR.n159 444.515
R2202 VDPWR.n274 VDPWR.n143 444.515
R2203 VDPWR.n265 VDPWR.n264 444.515
R2204 VDPWR.n251 VDPWR.n150 444.515
R2205 VDPWR.n604 VDPWR.n603 428.8
R2206 VDPWR.n357 VDPWR.n356 428.8
R2207 VDPWR.n421 VDPWR.n420 428.8
R2208 VDPWR.n247 VDPWR.n246 428.8
R2209 VDPWR.n275 VDPWR.n274 428.8
R2210 VDPWR.n264 VDPWR.n263 428.8
R2211 VDPWR.n252 VDPWR.n251 428.8
R2212 VDPWR.n603 VDPWR.n602 426.541
R2213 VDPWR.n356 VDPWR.n352 426.541
R2214 VDPWR.n422 VDPWR.n421 426.541
R2215 VDPWR.n246 VDPWR.n245 426.541
R2216 VDPWR.n276 VDPWR.n275 426.541
R2217 VDPWR.n263 VDPWR.n259 426.541
R2218 VDPWR.n253 VDPWR.n252 426.541
R2219 VDPWR.n616 VDPWR.n571 363.671
R2220 VDPWR.n443 VDPWR.n330 363.671
R2221 VDPWR.n415 VDPWR.n414 363.671
R2222 VDPWR.n198 VDPWR.n184 363.671
R2223 VDPWR.n112 VDPWR.n110 363.671
R2224 VDPWR.n125 VDPWR.n98 363.671
R2225 VDPWR.n181 VDPWR.n180 363.671
R2226 VDPWR.n629 VDPWR.n628 363.295
R2227 VDPWR.n456 VDPWR.n455 363.295
R2228 VDPWR.n413 VDPWR.n405 363.295
R2229 VDPWR.n224 VDPWR.n223 363.295
R2230 VDPWR.n277 VDPWR.n94 363.295
R2231 VDPWR.n319 VDPWR.n318 363.295
R2232 VDPWR.n227 VDPWR.n226 363.295
R2233 VDPWR.n616 VDPWR.n615 362.37
R2234 VDPWR.n415 VDPWR.n374 362.37
R2235 VDPWR.n443 VDPWR.n442 362.37
R2236 VDPWR.n199 VDPWR.n198 362.37
R2237 VDPWR.n180 VDPWR.n177 362.37
R2238 VDPWR.n118 VDPWR.n112 362.37
R2239 VDPWR.n127 VDPWR.n125 362.37
R2240 VDPWR.n628 VDPWR.n572 361.584
R2241 VDPWR.n405 VDPWR.n376 361.584
R2242 VDPWR.n455 VDPWR.n331 361.584
R2243 VDPWR.n223 VDPWR.n185 361.584
R2244 VDPWR.n228 VDPWR.n227 361.584
R2245 VDPWR.n278 VDPWR.n277 361.584
R2246 VDPWR.n318 VDPWR.n99 361.584
R2247 VDPWR.n626 VDPWR.n575 349.733
R2248 VDPWR.n403 VDPWR.n380 349.733
R2249 VDPWR.n453 VDPWR.n334 349.733
R2250 VDPWR.n619 VDPWR.n618 341.769
R2251 VDPWR.n417 VDPWR.n370 341.769
R2252 VDPWR.n446 VDPWR.n445 341.769
R2253 VDPWR.n428 VDPWR.n425 304.478
R2254 VDPWR.n580 VDPWR.n578 285.291
R2255 VDPWR.n401 VDPWR.n359 285.291
R2256 VDPWR.n339 VDPWR.n337 285.291
R2257 VDPWR.n607 VDPWR.n606 269.361
R2258 VDPWR.n371 VDPWR.n367 269.361
R2259 VDPWR.n427 VDPWR.n426 269.361
R2260 VDPWR.n684 VDPWR 190.871
R2261 VDPWR.n693 VDPWR 190.871
R2262 VDPWR.n684 VDPWR.n669 190.871
R2263 VDPWR.n700 VDPWR 190.871
R2264 VDPWR.n665 VDPWR 190.871
R2265 VDPWR.n700 VDPWR.n699 190.871
R2266 VDPWR VDPWR.n812 190.871
R2267 VDPWR.n812 VDPWR.n811 190.871
R2268 VDPWR VDPWR.n656 190.871
R2269 VDPWR.n828 VDPWR.n656 190.871
R2270 VDPWR.n786 VDPWR 190.871
R2271 VDPWR.n786 VDPWR.n785 190.871
R2272 VDPWR.n800 VDPWR 190.871
R2273 VDPWR.n800 VDPWR.n799 190.871
R2274 VDPWR.n760 VDPWR 190.871
R2275 VDPWR.n791 VDPWR 190.871
R2276 VDPWR.n760 VDPWR.n732 190.871
R2277 VDPWR.n752 VDPWR 190.871
R2278 VDPWR.n747 VDPWR 190.871
R2279 VDPWR.n752 VDPWR.n751 190.871
R2280 VDPWR.n688 VDPWR.n675 190.871
R2281 VDPWR VDPWR.n688 190.871
R2282 VDPWR.n689 VDPWR 190.871
R2283 VDPWR.n679 VDPWR.n678 190.871
R2284 VDPWR VDPWR.n679 190.871
R2285 VDPWR.n680 VDPWR 190.871
R2286 VDPWR.n725 VDPWR.n714 190.871
R2287 VDPWR VDPWR.n725 190.871
R2288 VDPWR.n721 VDPWR.n719 190.871
R2289 VDPWR VDPWR.n721 190.871
R2290 VDPWR.n764 VDPWR.n738 190.871
R2291 VDPWR VDPWR.n764 190.871
R2292 VDPWR.n765 VDPWR 190.871
R2293 VDPWR.n757 VDPWR 190.871
R2294 VDPWR VDPWR.n756 190.871
R2295 VDPWR.n756 VDPWR.n744 190.871
R2296 VDPWR.n504 VDPWR 190.871
R2297 VDPWR.n481 VDPWR 190.871
R2298 VDPWR.n504 VDPWR.n503 190.871
R2299 VDPWR.n477 VDPWR 190.871
R2300 VDPWR.n508 VDPWR 190.871
R2301 VDPWR.n477 VDPWR.n471 190.871
R2302 VDPWR.n487 VDPWR.n482 190.871
R2303 VDPWR.n487 VDPWR 190.871
R2304 VDPWR.n498 VDPWR 190.871
R2305 VDPWR.n494 VDPWR 190.871
R2306 VDPWR VDPWR.n493 190.871
R2307 VDPWR.n493 VDPWR.n492 190.871
R2308 VDPWR.n552 VDPWR 190.871
R2309 VDPWR.n529 VDPWR 190.871
R2310 VDPWR.n552 VDPWR.n551 190.871
R2311 VDPWR.n525 VDPWR 190.871
R2312 VDPWR.n556 VDPWR 190.871
R2313 VDPWR.n525 VDPWR.n519 190.871
R2314 VDPWR.n535 VDPWR.n530 190.871
R2315 VDPWR.n535 VDPWR 190.871
R2316 VDPWR.n546 VDPWR 190.871
R2317 VDPWR.n542 VDPWR 190.871
R2318 VDPWR VDPWR.n541 190.871
R2319 VDPWR.n541 VDPWR.n540 190.871
R2320 VDPWR.n603 VDPWR.n600 190.871
R2321 VDPWR.n600 VDPWR.n598 190.871
R2322 VDPWR.n355 VDPWR.n353 190.871
R2323 VDPWR.n356 VDPWR.n355 190.871
R2324 VDPWR.n396 VDPWR.n363 190.871
R2325 VDPWR.n421 VDPWR.n363 190.871
R2326 VDPWR.n7 VDPWR.n4 190.871
R2327 VDPWR.n7 VDPWR 190.871
R2328 VDPWR.n86 VDPWR 190.871
R2329 VDPWR.n77 VDPWR.n12 190.871
R2330 VDPWR VDPWR.n77 190.871
R2331 VDPWR.n78 VDPWR 190.871
R2332 VDPWR.n57 VDPWR.n26 190.871
R2333 VDPWR VDPWR.n26 190.871
R2334 VDPWR.n72 VDPWR.n16 190.871
R2335 VDPWR.n72 VDPWR 190.871
R2336 VDPWR.n49 VDPWR.n32 190.871
R2337 VDPWR VDPWR.n49 190.871
R2338 VDPWR.n50 VDPWR 190.871
R2339 VDPWR.n44 VDPWR 190.871
R2340 VDPWR VDPWR.n43 190.871
R2341 VDPWR.n43 VDPWR.n40 190.871
R2342 VDPWR.n246 VDPWR.n160 190.871
R2343 VDPWR.n217 VDPWR.n160 190.871
R2344 VDPWR.n275 VDPWR.n142 190.871
R2345 VDPWR.n142 VDPWR.n141 190.871
R2346 VDPWR.n262 VDPWR.n131 190.871
R2347 VDPWR.n263 VDPWR.n262 190.871
R2348 VDPWR.n237 VDPWR.n149 190.871
R2349 VDPWR.n252 VDPWR.n149 190.871
R2350 VDPWR.n694 VDPWR.n693 190.494
R2351 VDPWR.n698 VDPWR.n665 190.494
R2352 VDPWR.n792 VDPWR.n791 190.494
R2353 VDPWR.n750 VDPWR.n747 190.494
R2354 VDPWR.n689 VDPWR.n667 190.494
R2355 VDPWR.n680 VDPWR.n666 190.494
R2356 VDPWR.n765 VDPWR.n731 190.494
R2357 VDPWR.n757 VDPWR.n743 190.494
R2358 VDPWR.n502 VDPWR.n481 190.494
R2359 VDPWR.n509 VDPWR.n508 190.494
R2360 VDPWR.n499 VDPWR.n498 190.494
R2361 VDPWR.n494 VDPWR.n469 190.494
R2362 VDPWR.n550 VDPWR.n529 190.494
R2363 VDPWR.n557 VDPWR.n556 190.494
R2364 VDPWR.n547 VDPWR.n546 190.494
R2365 VDPWR.n542 VDPWR.n517 190.494
R2366 VDPWR.n87 VDPWR.n86 190.494
R2367 VDPWR.n78 VDPWR.n11 190.494
R2368 VDPWR.n50 VDPWR.n31 190.494
R2369 VDPWR.n44 VDPWR.n39 190.494
R2370 VDPWR.n46 VDPWR.n33 179.118
R2371 VDPWR.n47 VDPWR.n28 179.118
R2372 VDPWR.n52 VDPWR.n28 179.118
R2373 VDPWR.n55 VDPWR.n53 179.118
R2374 VDPWR.n55 VDPWR.n21 179.118
R2375 VDPWR.n69 VDPWR.n21 179.118
R2376 VDPWR.n69 VDPWR.n22 179.118
R2377 VDPWR.n22 VDPWR.n13 179.118
R2378 VDPWR.n74 VDPWR.n13 179.118
R2379 VDPWR.n75 VDPWR.n8 179.118
R2380 VDPWR.n80 VDPWR.n8 179.118
R2381 VDPWR.n81 VDPWR.n6 179.118
R2382 VDPWR.n213 VDPWR.n162 174.868
R2383 VDPWR.n316 VDPWR.n102 174.868
R2384 VDPWR.n42 VDPWR.n41 173.642
R2385 VDPWR.n85 VDPWR.n84 173.642
R2386 VDPWR.n214 VDPWR.n156 170.885
R2387 VDPWR.n308 VDPWR.n115 170.885
R2388 VDPWR.n267 VDPWR.n256 152.239
R2389 VDPWR.n242 VDPWR.n144 142.645
R2390 VDPWR.n281 VDPWR.n137 142.645
R2391 VDPWR.n581 VDPWR.n580 137.326
R2392 VDPWR.n340 VDPWR.n339 137.326
R2393 VDPWR.n608 VDPWR.n607 136.964
R2394 VDPWR.n371 VDPWR.n365 136.964
R2395 VDPWR.n201 VDPWR.n153 134.68
R2396 VDPWR.n302 VDPWR.n122 134.68
R2397 VDPWR.n824 VDPWR.n655 131.388
R2398 VDPWR.n829 VDPWR.n655 131.388
R2399 VDPWR.n809 VDPWR.n707 131.388
R2400 VDPWR.n810 VDPWR.n809 131.388
R2401 VDPWR.n778 VDPWR.n729 131.388
R2402 VDPWR.n798 VDPWR.n729 131.388
R2403 VDPWR.n783 VDPWR.n770 131.388
R2404 VDPWR.n784 VDPWR.n783 131.388
R2405 VDPWR.n718 VDPWR.n717 131.388
R2406 VDPWR.n722 VDPWR.n717 131.388
R2407 VDPWR.n819 VDPWR.n818 131.388
R2408 VDPWR.n818 VDPWR.n723 131.388
R2409 VDPWR.n61 VDPWR.n17 131.388
R2410 VDPWR.n71 VDPWR.n17 131.388
R2411 VDPWR.n60 VDPWR.n59 131.388
R2412 VDPWR.n59 VDPWR.n18 131.388
R2413 VDPWR.n425 VDPWR.n359 123.096
R2414 VDPWR.n428 VDPWR.n427 122.733
R2415 VDPWR.n75 VDPWR.n74 120.168
R2416 VDPWR.n47 VDPWR.n46 117.9
R2417 VDPWR.n81 VDPWR.n80 117.9
R2418 VDPWR VDPWR.n737 92.5005
R2419 VDPWR.n737 VDPWR.n735 92.5005
R2420 VDPWR.n738 VDPWR.n736 92.5005
R2421 VDPWR.n736 VDPWR.n735 92.5005
R2422 VDPWR VDPWR.n660 92.5005
R2423 VDPWR.n826 VDPWR.n660 92.5005
R2424 VDPWR VDPWR.n711 92.5005
R2425 VDPWR.n822 VDPWR.n711 92.5005
R2426 VDPWR.n815 VDPWR 92.5005
R2427 VDPWR.n815 VDPWR.n814 92.5005
R2428 VDPWR.n805 VDPWR.n714 92.5005
R2429 VDPWR.n814 VDPWR.n805 92.5005
R2430 VDPWR.n821 VDPWR.n820 92.5005
R2431 VDPWR.n822 VDPWR.n821 92.5005
R2432 VDPWR.n719 VDPWR.n704 92.5005
R2433 VDPWR.n826 VDPWR.n704 92.5005
R2434 VDPWR VDPWR.n677 92.5005
R2435 VDPWR.n677 VDPWR.n662 92.5005
R2436 VDPWR.n678 VDPWR.n676 92.5005
R2437 VDPWR.n676 VDPWR.n662 92.5005
R2438 VDPWR VDPWR.n674 92.5005
R2439 VDPWR.n674 VDPWR.n672 92.5005
R2440 VDPWR.n675 VDPWR.n673 92.5005
R2441 VDPWR.n673 VDPWR.n672 92.5005
R2442 VDPWR.n751 VDPWR.n746 92.5005
R2443 VDPWR.n746 VDPWR.n739 92.5005
R2444 VDPWR VDPWR.n745 92.5005
R2445 VDPWR.n745 VDPWR.n739 92.5005
R2446 VDPWR.n734 VDPWR.n732 92.5005
R2447 VDPWR.n735 VDPWR.n734 92.5005
R2448 VDPWR.n733 VDPWR 92.5005
R2449 VDPWR.n735 VDPWR.n733 92.5005
R2450 VDPWR.n799 VDPWR.n728 92.5005
R2451 VDPWR.n728 VDPWR.n726 92.5005
R2452 VDPWR.n773 VDPWR.n730 92.5005
R2453 VDPWR.n780 VDPWR.n773 92.5005
R2454 VDPWR.n785 VDPWR.n769 92.5005
R2455 VDPWR.n769 VDPWR.n767 92.5005
R2456 VDPWR VDPWR.n768 92.5005
R2457 VDPWR.n768 VDPWR.n767 92.5005
R2458 VDPWR.n779 VDPWR 92.5005
R2459 VDPWR.n780 VDPWR.n779 92.5005
R2460 VDPWR VDPWR.n727 92.5005
R2461 VDPWR.n727 VDPWR.n726 92.5005
R2462 VDPWR.n828 VDPWR.n827 92.5005
R2463 VDPWR.n827 VDPWR.n826 92.5005
R2464 VDPWR.n710 VDPWR.n654 92.5005
R2465 VDPWR.n822 VDPWR.n710 92.5005
R2466 VDPWR.n811 VDPWR.n804 92.5005
R2467 VDPWR.n814 VDPWR.n804 92.5005
R2468 VDPWR.n813 VDPWR 92.5005
R2469 VDPWR.n814 VDPWR.n813 92.5005
R2470 VDPWR VDPWR.n823 92.5005
R2471 VDPWR.n823 VDPWR.n822 92.5005
R2472 VDPWR.n825 VDPWR 92.5005
R2473 VDPWR.n826 VDPWR.n825 92.5005
R2474 VDPWR.n699 VDPWR.n664 92.5005
R2475 VDPWR.n664 VDPWR.n662 92.5005
R2476 VDPWR VDPWR.n663 92.5005
R2477 VDPWR.n663 VDPWR.n662 92.5005
R2478 VDPWR.n671 VDPWR.n669 92.5005
R2479 VDPWR.n672 VDPWR.n671 92.5005
R2480 VDPWR.n670 VDPWR 92.5005
R2481 VDPWR.n672 VDPWR.n670 92.5005
R2482 VDPWR VDPWR.n742 92.5005
R2483 VDPWR.n742 VDPWR.n739 92.5005
R2484 VDPWR.n744 VDPWR.n741 92.5005
R2485 VDPWR.n741 VDPWR.n739 92.5005
R2486 VDPWR.n484 VDPWR 92.5005
R2487 VDPWR.n489 VDPWR.n484 92.5005
R2488 VDPWR.n483 VDPWR.n482 92.5005
R2489 VDPWR.n485 VDPWR.n483 92.5005
R2490 VDPWR.n473 VDPWR.n471 92.5005
R2491 VDPWR.n476 VDPWR.n473 92.5005
R2492 VDPWR.n472 VDPWR 92.5005
R2493 VDPWR.n474 VDPWR.n472 92.5005
R2494 VDPWR.n503 VDPWR.n480 92.5005
R2495 VDPWR.n480 VDPWR.n476 92.5005
R2496 VDPWR VDPWR.n479 92.5005
R2497 VDPWR.n479 VDPWR.n474 92.5005
R2498 VDPWR VDPWR.n491 92.5005
R2499 VDPWR.n491 VDPWR.n489 92.5005
R2500 VDPWR.n492 VDPWR.n490 92.5005
R2501 VDPWR.n490 VDPWR.n485 92.5005
R2502 VDPWR.n532 VDPWR 92.5005
R2503 VDPWR.n537 VDPWR.n532 92.5005
R2504 VDPWR.n531 VDPWR.n530 92.5005
R2505 VDPWR.n533 VDPWR.n531 92.5005
R2506 VDPWR.n521 VDPWR.n519 92.5005
R2507 VDPWR.n524 VDPWR.n521 92.5005
R2508 VDPWR.n520 VDPWR 92.5005
R2509 VDPWR.n522 VDPWR.n520 92.5005
R2510 VDPWR.n551 VDPWR.n528 92.5005
R2511 VDPWR.n528 VDPWR.n524 92.5005
R2512 VDPWR VDPWR.n527 92.5005
R2513 VDPWR.n527 VDPWR.n522 92.5005
R2514 VDPWR VDPWR.n539 92.5005
R2515 VDPWR.n539 VDPWR.n537 92.5005
R2516 VDPWR.n540 VDPWR.n538 92.5005
R2517 VDPWR.n538 VDPWR.n533 92.5005
R2518 VDPWR VDPWR.n30 92.5005
R2519 VDPWR.n30 VDPWR.n28 92.5005
R2520 VDPWR.n32 VDPWR.n29 92.5005
R2521 VDPWR.n29 VDPWR.n28 92.5005
R2522 VDPWR VDPWR.n15 92.5005
R2523 VDPWR.n15 VDPWR.n13 92.5005
R2524 VDPWR VDPWR.n70 92.5005
R2525 VDPWR.n70 VDPWR.n69 92.5005
R2526 VDPWR.n54 VDPWR 92.5005
R2527 VDPWR.n55 VDPWR.n54 92.5005
R2528 VDPWR.n57 VDPWR.n56 92.5005
R2529 VDPWR.n56 VDPWR.n55 92.5005
R2530 VDPWR.n68 VDPWR.n67 92.5005
R2531 VDPWR.n69 VDPWR.n68 92.5005
R2532 VDPWR.n16 VDPWR.n14 92.5005
R2533 VDPWR.n14 VDPWR.n13 92.5005
R2534 VDPWR VDPWR.n10 92.5005
R2535 VDPWR.n10 VDPWR.n8 92.5005
R2536 VDPWR.n12 VDPWR.n9 92.5005
R2537 VDPWR.n9 VDPWR.n8 92.5005
R2538 VDPWR.n83 VDPWR 92.5005
R2539 VDPWR.n5 VDPWR.n4 92.5005
R2540 VDPWR.n6 VDPWR.n5 92.5005
R2541 VDPWR VDPWR.n35 92.5005
R2542 VDPWR.n35 VDPWR.n33 92.5005
R2543 VDPWR.n40 VDPWR.n34 92.5005
R2544 VDPWR.n506 VDPWR.n474 91.6935
R2545 VDPWR.n506 VDPWR.n476 91.6935
R2546 VDPWR.n496 VDPWR.n485 91.6935
R2547 VDPWR.n496 VDPWR.n489 91.6935
R2548 VDPWR.n554 VDPWR.n522 91.6935
R2549 VDPWR.n554 VDPWR.n524 91.6935
R2550 VDPWR.n544 VDPWR.n533 91.6935
R2551 VDPWR.n544 VDPWR.n537 91.6935
R2552 VDPWR.n754 VDPWR.n739 89.559
R2553 VDPWR.n759 VDPWR.n739 89.559
R2554 VDPWR.n762 VDPWR.n735 89.559
R2555 VDPWR.n789 VDPWR.n735 89.559
R2556 VDPWR.n788 VDPWR.n767 89.559
R2557 VDPWR.n781 VDPWR.n767 89.559
R2558 VDPWR.n781 VDPWR.n780 89.559
R2559 VDPWR.n780 VDPWR.n774 89.559
R2560 VDPWR.n774 VDPWR.n726 89.559
R2561 VDPWR.n802 VDPWR.n726 89.559
R2562 VDPWR.n814 VDPWR.n803 89.559
R2563 VDPWR.n814 VDPWR.n709 89.559
R2564 VDPWR.n822 VDPWR.n709 89.559
R2565 VDPWR.n822 VDPWR.n659 89.559
R2566 VDPWR.n826 VDPWR.n659 89.559
R2567 VDPWR.n826 VDPWR.n703 89.559
R2568 VDPWR.n702 VDPWR.n662 89.559
R2569 VDPWR.n683 VDPWR.n662 89.559
R2570 VDPWR.n686 VDPWR.n672 89.559
R2571 VDPWR.n691 VDPWR.n672 89.559
R2572 VDPWR.n590 VDPWR.n589 85.0829
R2573 VDPWR.n590 VDPWR.n571 85.0829
R2574 VDPWR.n435 VDPWR.n330 85.0829
R2575 VDPWR.n436 VDPWR.n435 85.0829
R2576 VDPWR.n414 VDPWR.n375 85.0829
R2577 VDPWR.n390 VDPWR.n375 85.0829
R2578 VDPWR.n209 VDPWR.n188 85.0829
R2579 VDPWR.n209 VDPWR.n184 85.0829
R2580 VDPWR.n313 VDPWR.n312 85.0829
R2581 VDPWR.n312 VDPWR.n110 85.0829
R2582 VDPWR.n295 VDPWR.n98 85.0829
R2583 VDPWR.n296 VDPWR.n295 85.0829
R2584 VDPWR.n181 VDPWR.n175 85.0829
R2585 VDPWR.n175 VDPWR.n174 85.0829
R2586 VDPWR.n84 VDPWR.n83 79.4196
R2587 VDPWR.n41 VDPWR.n34 79.4196
R2588 VDPWR.n598 VDPWR.n582 66.7857
R2589 VDPWR.n353 VDPWR.n341 66.7857
R2590 VDPWR.n397 VDPWR.n396 66.7857
R2591 VDPWR.n218 VDPWR.n217 66.7857
R2592 VDPWR.n141 VDPWR.n108 66.7857
R2593 VDPWR.n291 VDPWR.n131 66.7857
R2594 VDPWR.n238 VDPWR.n237 66.7857
R2595 VDPWR.n610 VDPWR.n596 66.1931
R2596 VDPWR.n431 VDPWR.n345 66.1931
R2597 VDPWR.n395 VDPWR.n394 66.1931
R2598 VDPWR.n216 VDPWR.n192 66.1931
R2599 VDPWR.n140 VDPWR.n117 66.1931
R2600 VDPWR.n130 VDPWR.n129 66.1931
R2601 VDPWR.n236 VDPWR.n235 66.1931
R2602 VDPWR.n618 VDPWR.n587 62.6339
R2603 VDPWR.n418 VDPWR.n417 62.6339
R2604 VDPWR.n445 VDPWR.n346 62.6339
R2605 VDPWR.n256 VDPWR.n144 61.5478
R2606 VDPWR.n287 VDPWR.n137 61.5478
R2607 VDPWR.n201 VDPWR.n200 61.3667
R2608 VDPWR.n267 VDPWR.n122 61.3667
R2609 VDPWR.n626 VDPWR.n625 60.4616
R2610 VDPWR.n403 VDPWR.n402 60.4616
R2611 VDPWR.n453 VDPWR.n452 60.4616
R2612 VDPWR.n789 VDPWR.n788 60.084
R2613 VDPWR.n803 VDPWR.n802 60.084
R2614 VDPWR.n703 VDPWR.n702 60.084
R2615 VDPWR VDPWR.n707 59.4829
R2616 VDPWR VDPWR.n707 59.4829
R2617 VDPWR.n824 VDPWR 59.4829
R2618 VDPWR VDPWR.n824 59.4829
R2619 VDPWR.n811 VDPWR.n810 59.4829
R2620 VDPWR.n810 VDPWR.n654 59.4829
R2621 VDPWR.n829 VDPWR.n828 59.4829
R2622 VDPWR.n770 VDPWR 59.4829
R2623 VDPWR VDPWR.n770 59.4829
R2624 VDPWR VDPWR.n778 59.4829
R2625 VDPWR.n778 VDPWR 59.4829
R2626 VDPWR.n785 VDPWR.n784 59.4829
R2627 VDPWR.n784 VDPWR.n730 59.4829
R2628 VDPWR.n799 VDPWR.n798 59.4829
R2629 VDPWR.n819 VDPWR.n714 59.4829
R2630 VDPWR.n820 VDPWR.n819 59.4829
R2631 VDPWR.n719 VDPWR.n718 59.4829
R2632 VDPWR VDPWR.n723 59.4829
R2633 VDPWR.n723 VDPWR 59.4829
R2634 VDPWR VDPWR.n722 59.4829
R2635 VDPWR.n722 VDPWR 59.4829
R2636 VDPWR.n60 VDPWR.n57 59.4829
R2637 VDPWR.n67 VDPWR.n60 59.4829
R2638 VDPWR.n61 VDPWR.n16 59.4829
R2639 VDPWR VDPWR.n18 59.4829
R2640 VDPWR VDPWR.n18 59.4829
R2641 VDPWR.n71 VDPWR 59.4829
R2642 VDPWR VDPWR.n71 59.4829
R2643 VDPWR.n830 VDPWR.n829 59.1064
R2644 VDPWR.n798 VDPWR.n797 59.1064
R2645 VDPWR.n718 VDPWR.n652 59.1064
R2646 VDPWR.n66 VDPWR.n61 59.1064
R2647 VDPWR.n762 VDPWR.n759 58.9504
R2648 VDPWR.n686 VDPWR.n683 58.9504
R2649 VDPWR.n589 VDPWR.n588 52.3937
R2650 VDPWR.n436 VDPWR.n432 52.3937
R2651 VDPWR.n390 VDPWR.n386 52.3937
R2652 VDPWR.n219 VDPWR.n188 52.3937
R2653 VDPWR.n314 VDPWR.n313 52.3937
R2654 VDPWR.n296 VDPWR.n292 52.3937
R2655 VDPWR.n174 VDPWR.n167 52.3937
R2656 VDPWR.n611 VDPWR.n586 51.2005
R2657 VDPWR.n438 VDPWR.n437 51.2005
R2658 VDPWR.n392 VDPWR.n391 51.2005
R2659 VDPWR.n205 VDPWR.n204 51.2005
R2660 VDPWR.n306 VDPWR.n109 51.2005
R2661 VDPWR.n298 VDPWR.n297 51.2005
R2662 VDPWR.n233 VDPWR.n170 51.2005
R2663 VDPWR.n622 VDPWR.n621 37.0005
R2664 VDPWR.n621 VDPWR.n578 37.0005
R2665 VDPWR.n574 VDPWR.n572 37.0005
R2666 VDPWR.n580 VDPWR.n574 37.0005
R2667 VDPWR.n615 VDPWR.n594 37.0005
R2668 VDPWR.n607 VDPWR.n594 37.0005
R2669 VDPWR.n613 VDPWR.n585 37.0005
R2670 VDPWR.n606 VDPWR.n585 37.0005
R2671 VDPWR.n591 VDPWR.n590 37.0005
R2672 VDPWR.n591 VDPWR.n575 37.0005
R2673 VDPWR.n449 VDPWR.n448 37.0005
R2674 VDPWR.n448 VDPWR.n337 37.0005
R2675 VDPWR.n440 VDPWR.n344 37.0005
R2676 VDPWR.n426 VDPWR.n344 37.0005
R2677 VDPWR.n377 VDPWR.n376 37.0005
R2678 VDPWR.n377 VDPWR.n359 37.0005
R2679 VDPWR.n374 VDPWR.n372 37.0005
R2680 VDPWR.n372 VDPWR.n371 37.0005
R2681 VDPWR.n435 VDPWR.n434 37.0005
R2682 VDPWR.n434 VDPWR.n334 37.0005
R2683 VDPWR.n333 VDPWR.n331 37.0005
R2684 VDPWR.n339 VDPWR.n333 37.0005
R2685 VDPWR.n442 VDPWR.n348 37.0005
R2686 VDPWR.n427 VDPWR.n348 37.0005
R2687 VDPWR.n400 VDPWR.n399 37.0005
R2688 VDPWR.n401 VDPWR.n400 37.0005
R2689 VDPWR.n389 VDPWR.n388 37.0005
R2690 VDPWR.n388 VDPWR.n367 37.0005
R2691 VDPWR.n381 VDPWR.n375 37.0005
R2692 VDPWR.n381 VDPWR.n380 37.0005
R2693 VDPWR.n280 VDPWR.n132 37.0005
R2694 VDPWR.n281 VDPWR.n280 37.0005
R2695 VDPWR.n301 VDPWR.n300 37.0005
R2696 VDPWR.n302 VDPWR.n301 37.0005
R2697 VDPWR.n229 VDPWR.n228 37.0005
R2698 VDPWR.n229 VDPWR.n144 37.0005
R2699 VDPWR.n177 VDPWR.n171 37.0005
R2700 VDPWR.n201 VDPWR.n171 37.0005
R2701 VDPWR.n295 VDPWR.n294 37.0005
R2702 VDPWR.n294 VDPWR.n102 37.0005
R2703 VDPWR.n101 VDPWR.n99 37.0005
R2704 VDPWR.n137 VDPWR.n101 37.0005
R2705 VDPWR.n127 VDPWR.n126 37.0005
R2706 VDPWR.n126 VDPWR.n122 37.0005
R2707 VDPWR.n210 VDPWR.n209 37.0005
R2708 VDPWR.n213 VDPWR.n210 37.0005
R2709 VDPWR.n221 VDPWR.n185 37.0005
R2710 VDPWR.n221 VDPWR.n144 37.0005
R2711 VDPWR.n202 VDPWR.n199 37.0005
R2712 VDPWR.n202 VDPWR.n201 37.0005
R2713 VDPWR.n312 VDPWR.n311 37.0005
R2714 VDPWR.n311 VDPWR.n102 37.0005
R2715 VDPWR.n278 VDPWR.n107 37.0005
R2716 VDPWR.n137 VDPWR.n107 37.0005
R2717 VDPWR.n118 VDPWR.n111 37.0005
R2718 VDPWR.n122 VDPWR.n111 37.0005
R2719 VDPWR.n190 VDPWR.n164 37.0005
R2720 VDPWR.n242 VDPWR.n164 37.0005
R2721 VDPWR.n196 VDPWR.n193 37.0005
R2722 VDPWR.n193 VDPWR.n153 37.0005
R2723 VDPWR.n283 VDPWR.n282 37.0005
R2724 VDPWR.n282 VDPWR.n281 37.0005
R2725 VDPWR.n304 VDPWR.n303 37.0005
R2726 VDPWR.n303 VDPWR.n302 37.0005
R2727 VDPWR.n241 VDPWR.n240 37.0005
R2728 VDPWR.n242 VDPWR.n241 37.0005
R2729 VDPWR.n169 VDPWR.n168 37.0005
R2730 VDPWR.n168 VDPWR.n153 37.0005
R2731 VDPWR.n175 VDPWR.n172 37.0005
R2732 VDPWR.n213 VDPWR.n172 37.0005
R2733 VDPWR.n249 VDPWR.n156 31.3172
R2734 VDPWR.n308 VDPWR.n113 31.3172
R2735 VDPWR.n243 VDPWR.n162 30.2311
R2736 VDPWR.n316 VDPWR.n105 30.2311
R2737 VDPWR.n614 VDPWR.n595 26.6787
R2738 VDPWR.n441 VDPWR.n349 26.6787
R2739 VDPWR.n387 VDPWR.n364 26.6787
R2740 VDPWR.n197 VDPWR.n159 26.6787
R2741 VDPWR.n143 VDPWR.n119 26.6787
R2742 VDPWR.n265 VDPWR.n128 26.6787
R2743 VDPWR.n176 VDPWR.n150 26.6787
R2744 VDPWR.n601 VDPWR.n583 26.63
R2745 VDPWR.n351 VDPWR.n342 26.63
R2746 VDPWR.n423 VDPWR.n362 26.63
R2747 VDPWR.n189 VDPWR.n161 26.63
R2748 VDPWR.n285 VDPWR.n284 26.63
R2749 VDPWR.n136 VDPWR.n135 26.63
R2750 VDPWR.n254 VDPWR.n148 26.63
R2751 VDPWR.n485 VDPWR.n476 26.5564
R2752 VDPWR.n533 VDPWR.n524 26.5564
R2753 VDPWR.n766 VDPWR.n765 23.1255
R2754 VDPWR.n789 VDPWR.n766 23.1255
R2755 VDPWR.n764 VDPWR.n763 23.1255
R2756 VDPWR.n763 VDPWR.n762 23.1255
R2757 VDPWR.n818 VDPWR.n817 23.1255
R2758 VDPWR.n817 VDPWR.n709 23.1255
R2759 VDPWR.n717 VDPWR.n716 23.1255
R2760 VDPWR.n716 VDPWR.n659 23.1255
R2761 VDPWR.n721 VDPWR.n720 23.1255
R2762 VDPWR.n720 VDPWR.n703 23.1255
R2763 VDPWR.n725 VDPWR.n724 23.1255
R2764 VDPWR.n803 VDPWR.n724 23.1255
R2765 VDPWR.n681 VDPWR.n680 23.1255
R2766 VDPWR.n683 VDPWR.n681 23.1255
R2767 VDPWR.n679 VDPWR.n661 23.1255
R2768 VDPWR.n702 VDPWR.n661 23.1255
R2769 VDPWR.n690 VDPWR.n689 23.1255
R2770 VDPWR.n691 VDPWR.n690 23.1255
R2771 VDPWR.n688 VDPWR.n687 23.1255
R2772 VDPWR.n687 VDPWR.n686 23.1255
R2773 VDPWR.n747 VDPWR.n740 23.1255
R2774 VDPWR.n759 VDPWR.n740 23.1255
R2775 VDPWR.n753 VDPWR.n752 23.1255
R2776 VDPWR.n754 VDPWR.n753 23.1255
R2777 VDPWR.n791 VDPWR.n790 23.1255
R2778 VDPWR.n790 VDPWR.n789 23.1255
R2779 VDPWR.n761 VDPWR.n760 23.1255
R2780 VDPWR.n762 VDPWR.n761 23.1255
R2781 VDPWR.n783 VDPWR.n782 23.1255
R2782 VDPWR.n782 VDPWR.n781 23.1255
R2783 VDPWR.n776 VDPWR.n729 23.1255
R2784 VDPWR.n776 VDPWR.n774 23.1255
R2785 VDPWR.n801 VDPWR.n800 23.1255
R2786 VDPWR.n802 VDPWR.n801 23.1255
R2787 VDPWR.n787 VDPWR.n786 23.1255
R2788 VDPWR.n788 VDPWR.n787 23.1255
R2789 VDPWR.n809 VDPWR.n808 23.1255
R2790 VDPWR.n808 VDPWR.n709 23.1255
R2791 VDPWR.n705 VDPWR.n655 23.1255
R2792 VDPWR.n705 VDPWR.n659 23.1255
R2793 VDPWR.n658 VDPWR.n656 23.1255
R2794 VDPWR.n703 VDPWR.n658 23.1255
R2795 VDPWR.n812 VDPWR.n806 23.1255
R2796 VDPWR.n806 VDPWR.n803 23.1255
R2797 VDPWR.n682 VDPWR.n665 23.1255
R2798 VDPWR.n683 VDPWR.n682 23.1255
R2799 VDPWR.n701 VDPWR.n700 23.1255
R2800 VDPWR.n702 VDPWR.n701 23.1255
R2801 VDPWR.n693 VDPWR.n692 23.1255
R2802 VDPWR.n692 VDPWR.n691 23.1255
R2803 VDPWR.n685 VDPWR.n684 23.1255
R2804 VDPWR.n686 VDPWR.n685 23.1255
R2805 VDPWR.n758 VDPWR.n757 23.1255
R2806 VDPWR.n759 VDPWR.n758 23.1255
R2807 VDPWR.n756 VDPWR.n755 23.1255
R2808 VDPWR.n755 VDPWR.n754 23.1255
R2809 VDPWR.n498 VDPWR.n497 23.1255
R2810 VDPWR.n497 VDPWR.n496 23.1255
R2811 VDPWR.n488 VDPWR.n487 23.1255
R2812 VDPWR.n496 VDPWR.n488 23.1255
R2813 VDPWR.n508 VDPWR.n507 23.1255
R2814 VDPWR.n507 VDPWR.n506 23.1255
R2815 VDPWR.n478 VDPWR.n477 23.1255
R2816 VDPWR.n506 VDPWR.n478 23.1255
R2817 VDPWR.n481 VDPWR.n475 23.1255
R2818 VDPWR.n506 VDPWR.n475 23.1255
R2819 VDPWR.n505 VDPWR.n504 23.1255
R2820 VDPWR.n506 VDPWR.n505 23.1255
R2821 VDPWR.n495 VDPWR.n494 23.1255
R2822 VDPWR.n496 VDPWR.n495 23.1255
R2823 VDPWR.n493 VDPWR.n486 23.1255
R2824 VDPWR.n496 VDPWR.n486 23.1255
R2825 VDPWR.n546 VDPWR.n545 23.1255
R2826 VDPWR.n545 VDPWR.n544 23.1255
R2827 VDPWR.n536 VDPWR.n535 23.1255
R2828 VDPWR.n544 VDPWR.n536 23.1255
R2829 VDPWR.n556 VDPWR.n555 23.1255
R2830 VDPWR.n555 VDPWR.n554 23.1255
R2831 VDPWR.n526 VDPWR.n525 23.1255
R2832 VDPWR.n554 VDPWR.n526 23.1255
R2833 VDPWR.n529 VDPWR.n523 23.1255
R2834 VDPWR.n554 VDPWR.n523 23.1255
R2835 VDPWR.n553 VDPWR.n552 23.1255
R2836 VDPWR.n554 VDPWR.n553 23.1255
R2837 VDPWR.n543 VDPWR.n542 23.1255
R2838 VDPWR.n544 VDPWR.n543 23.1255
R2839 VDPWR.n541 VDPWR.n534 23.1255
R2840 VDPWR.n544 VDPWR.n534 23.1255
R2841 VDPWR.n51 VDPWR.n50 23.1255
R2842 VDPWR.n52 VDPWR.n51 23.1255
R2843 VDPWR.n49 VDPWR.n48 23.1255
R2844 VDPWR.n48 VDPWR.n47 23.1255
R2845 VDPWR.n59 VDPWR.n58 23.1255
R2846 VDPWR.n58 VDPWR.n21 23.1255
R2847 VDPWR.n24 VDPWR.n17 23.1255
R2848 VDPWR.n24 VDPWR.n22 23.1255
R2849 VDPWR.n73 VDPWR.n72 23.1255
R2850 VDPWR.n74 VDPWR.n73 23.1255
R2851 VDPWR.n27 VDPWR.n26 23.1255
R2852 VDPWR.n53 VDPWR.n27 23.1255
R2853 VDPWR.n79 VDPWR.n78 23.1255
R2854 VDPWR.n80 VDPWR.n79 23.1255
R2855 VDPWR.n77 VDPWR.n76 23.1255
R2856 VDPWR.n76 VDPWR.n75 23.1255
R2857 VDPWR.n86 VDPWR.n85 23.1255
R2858 VDPWR.n82 VDPWR.n7 23.1255
R2859 VDPWR.n82 VDPWR.n81 23.1255
R2860 VDPWR.n45 VDPWR.n44 23.1255
R2861 VDPWR.n46 VDPWR.n45 23.1255
R2862 VDPWR.n43 VDPWR.n42 23.1255
R2863 VDPWR.n612 VDPWR.n611 19.0689
R2864 VDPWR.n439 VDPWR.n438 19.0689
R2865 VDPWR.n393 VDPWR.n392 19.0689
R2866 VDPWR.n204 VDPWR.n194 19.0689
R2867 VDPWR.n306 VDPWR.n305 19.0689
R2868 VDPWR.n299 VDPWR.n298 19.0689
R2869 VDPWR.n234 VDPWR.n233 19.0689
R2870 VDPWR.n606 VDPWR.n587 17.7406
R2871 VDPWR.n418 VDPWR.n367 17.7406
R2872 VDPWR.n426 VDPWR.n346 17.7406
R2873 VDPWR.n622 VDPWR.n583 17.4344
R2874 VDPWR.n449 VDPWR.n342 17.4344
R2875 VDPWR.n399 VDPWR.n362 17.4344
R2876 VDPWR.n190 VDPWR.n189 17.4344
R2877 VDPWR.n284 VDPWR.n283 17.4344
R2878 VDPWR.n135 VDPWR.n132 17.4344
R2879 VDPWR.n240 VDPWR.n148 17.4344
R2880 VDPWR.n588 VDPWR.n582 16.8923
R2881 VDPWR.n397 VDPWR.n386 16.8923
R2882 VDPWR.n432 VDPWR.n341 16.8923
R2883 VDPWR.n238 VDPWR.n167 16.8923
R2884 VDPWR.n219 VDPWR.n218 16.8923
R2885 VDPWR.n314 VDPWR.n108 16.8923
R2886 VDPWR.n292 VDPWR.n291 16.8923
R2887 VDPWR.n614 VDPWR.n613 16.6793
R2888 VDPWR.n441 VDPWR.n440 16.6793
R2889 VDPWR.n389 VDPWR.n387 16.6793
R2890 VDPWR.n197 VDPWR.n196 16.6793
R2891 VDPWR.n304 VDPWR.n119 16.6793
R2892 VDPWR.n300 VDPWR.n128 16.6793
R2893 VDPWR.n176 VDPWR.n169 16.6793
R2894 VDPWR.n608 VDPWR.n595 14.2313
R2895 VDPWR.n600 VDPWR.n599 14.2313
R2896 VDPWR.n599 VDPWR.n575 14.2313
R2897 VDPWR.n601 VDPWR.n581 14.2313
R2898 VDPWR.n355 VDPWR.n354 14.2313
R2899 VDPWR.n354 VDPWR.n334 14.2313
R2900 VDPWR.n351 VDPWR.n340 14.2313
R2901 VDPWR.n429 VDPWR.n349 14.2313
R2902 VDPWR.n429 VDPWR.n428 14.2313
R2903 VDPWR.n424 VDPWR.n423 14.2313
R2904 VDPWR.n425 VDPWR.n424 14.2313
R2905 VDPWR.n379 VDPWR.n363 14.2313
R2906 VDPWR.n380 VDPWR.n379 14.2313
R2907 VDPWR.n365 VDPWR.n364 14.2313
R2908 VDPWR.n262 VDPWR.n261 14.2313
R2909 VDPWR.n261 VDPWR.n102 14.2313
R2910 VDPWR.n288 VDPWR.n136 14.2313
R2911 VDPWR.n288 VDPWR.n287 14.2313
R2912 VDPWR.n266 VDPWR.n265 14.2313
R2913 VDPWR.n267 VDPWR.n266 14.2313
R2914 VDPWR.n212 VDPWR.n160 14.2313
R2915 VDPWR.n213 VDPWR.n212 14.2313
R2916 VDPWR.n161 VDPWR.n145 14.2313
R2917 VDPWR.n256 VDPWR.n145 14.2313
R2918 VDPWR.n159 VDPWR.n157 14.2313
R2919 VDPWR.n200 VDPWR.n157 14.2313
R2920 VDPWR.n271 VDPWR.n142 14.2313
R2921 VDPWR.n271 VDPWR.n102 14.2313
R2922 VDPWR.n286 VDPWR.n285 14.2313
R2923 VDPWR.n287 VDPWR.n286 14.2313
R2924 VDPWR.n268 VDPWR.n143 14.2313
R2925 VDPWR.n268 VDPWR.n267 14.2313
R2926 VDPWR.n255 VDPWR.n254 14.2313
R2927 VDPWR.n256 VDPWR.n255 14.2313
R2928 VDPWR.n208 VDPWR.n149 14.2313
R2929 VDPWR.n213 VDPWR.n208 14.2313
R2930 VDPWR.n151 VDPWR.n150 14.2313
R2931 VDPWR.n200 VDPWR.n151 14.2313
R2932 VDPWR.n84 VDPWR.n6 8.97701
R2933 VDPWR.n41 VDPWR.n33 8.97701
R2934 VDPWR.n249 VDPWR.n153 8.87055
R2935 VDPWR.n302 VDPWR.n113 8.87055
R2936 VDPWR.n619 VDPWR.n575 7.96544
R2937 VDPWR.n380 VDPWR.n370 7.96544
R2938 VDPWR.n446 VDPWR.n334 7.96544
R2939 VDPWR.n611 VDPWR.n593 7.11588
R2940 VDPWR.n618 VDPWR.n593 7.11588
R2941 VDPWR.n588 VDPWR.n576 7.11588
R2942 VDPWR.n626 VDPWR.n576 7.11588
R2943 VDPWR.n628 VDPWR.n627 7.11588
R2944 VDPWR.n627 VDPWR.n626 7.11588
R2945 VDPWR.n617 VDPWR.n616 7.11588
R2946 VDPWR.n618 VDPWR.n617 7.11588
R2947 VDPWR.n432 VDPWR.n335 7.11588
R2948 VDPWR.n453 VDPWR.n335 7.11588
R2949 VDPWR.n438 VDPWR.n347 7.11588
R2950 VDPWR.n445 VDPWR.n347 7.11588
R2951 VDPWR.n444 VDPWR.n443 7.11588
R2952 VDPWR.n445 VDPWR.n444 7.11588
R2953 VDPWR.n455 VDPWR.n454 7.11588
R2954 VDPWR.n454 VDPWR.n453 7.11588
R2955 VDPWR.n386 VDPWR.n383 7.11588
R2956 VDPWR.n403 VDPWR.n383 7.11588
R2957 VDPWR.n392 VDPWR.n369 7.11588
R2958 VDPWR.n417 VDPWR.n369 7.11588
R2959 VDPWR.n416 VDPWR.n415 7.11588
R2960 VDPWR.n417 VDPWR.n416 7.11588
R2961 VDPWR.n405 VDPWR.n404 7.11588
R2962 VDPWR.n404 VDPWR.n403 7.11588
R2963 VDPWR.n292 VDPWR.n104 7.11588
R2964 VDPWR.n316 VDPWR.n104 7.11588
R2965 VDPWR.n298 VDPWR.n114 7.11588
R2966 VDPWR.n308 VDPWR.n114 7.11588
R2967 VDPWR.n125 VDPWR.n116 7.11588
R2968 VDPWR.n308 VDPWR.n116 7.11588
R2969 VDPWR.n318 VDPWR.n317 7.11588
R2970 VDPWR.n317 VDPWR.n316 7.11588
R2971 VDPWR.n223 VDPWR.n222 7.11588
R2972 VDPWR.n222 VDPWR.n162 7.11588
R2973 VDPWR.n198 VDPWR.n195 7.11588
R2974 VDPWR.n195 VDPWR.n156 7.11588
R2975 VDPWR.n204 VDPWR.n203 7.11588
R2976 VDPWR.n203 VDPWR.n156 7.11588
R2977 VDPWR.n220 VDPWR.n219 7.11588
R2978 VDPWR.n220 VDPWR.n162 7.11588
R2979 VDPWR.n277 VDPWR.n103 7.11588
R2980 VDPWR.n316 VDPWR.n103 7.11588
R2981 VDPWR.n309 VDPWR.n112 7.11588
R2982 VDPWR.n309 VDPWR.n308 7.11588
R2983 VDPWR.n307 VDPWR.n306 7.11588
R2984 VDPWR.n308 VDPWR.n307 7.11588
R2985 VDPWR.n315 VDPWR.n314 7.11588
R2986 VDPWR.n316 VDPWR.n315 7.11588
R2987 VDPWR.n230 VDPWR.n167 7.11588
R2988 VDPWR.n230 VDPWR.n162 7.11588
R2989 VDPWR.n233 VDPWR.n232 7.11588
R2990 VDPWR.n232 VDPWR.n156 7.11588
R2991 VDPWR.n180 VDPWR.n179 7.11588
R2992 VDPWR.n179 VDPWR.n156 7.11588
R2993 VDPWR.n227 VDPWR.n173 7.11588
R2994 VDPWR.n173 VDPWR.n162 7.11588
R2995 VDPWR.n323 VDPWR 6.74008
R2996 VDPWR.n460 VDPWR 6.737
R2997 VDPWR.n323 VDPWR 6.73352
R2998 VDPWR.n409 VDPWR.n408 6.63939
R2999 VDPWR.n634 VDPWR.n633 6.63939
R3000 VDPWR.n596 VDPWR.n584 5.78175
R3001 VDPWR.n619 VDPWR.n584 5.78175
R3002 VDPWR.n610 VDPWR.n609 5.78175
R3003 VDPWR.n609 VDPWR.n587 5.78175
R3004 VDPWR.n605 VDPWR.n604 5.78175
R3005 VDPWR.n605 VDPWR.n587 5.78175
R3006 VDPWR.n602 VDPWR.n577 5.78175
R3007 VDPWR.n625 VDPWR.n577 5.78175
R3008 VDPWR.n624 VDPWR.n623 5.78175
R3009 VDPWR.n625 VDPWR.n624 5.78175
R3010 VDPWR.n620 VDPWR.n586 5.78175
R3011 VDPWR.n620 VDPWR.n619 5.78175
R3012 VDPWR.n352 VDPWR.n336 5.78175
R3013 VDPWR.n452 VDPWR.n336 5.78175
R3014 VDPWR.n358 VDPWR.n357 5.78175
R3015 VDPWR.n358 VDPWR.n346 5.78175
R3016 VDPWR.n431 VDPWR.n430 5.78175
R3017 VDPWR.n430 VDPWR.n346 5.78175
R3018 VDPWR.n451 VDPWR.n450 5.78175
R3019 VDPWR.n452 VDPWR.n451 5.78175
R3020 VDPWR.n447 VDPWR.n345 5.78175
R3021 VDPWR.n447 VDPWR.n446 5.78175
R3022 VDPWR.n437 VDPWR.n343 5.78175
R3023 VDPWR.n446 VDPWR.n343 5.78175
R3024 VDPWR.n398 VDPWR.n360 5.78175
R3025 VDPWR.n402 VDPWR.n360 5.78175
R3026 VDPWR.n394 VDPWR.n368 5.78175
R3027 VDPWR.n418 VDPWR.n368 5.78175
R3028 VDPWR.n395 VDPWR.n385 5.78175
R3029 VDPWR.n385 VDPWR.n370 5.78175
R3030 VDPWR.n422 VDPWR.n361 5.78175
R3031 VDPWR.n402 VDPWR.n361 5.78175
R3032 VDPWR.n420 VDPWR.n419 5.78175
R3033 VDPWR.n419 VDPWR.n418 5.78175
R3034 VDPWR.n391 VDPWR.n384 5.78175
R3035 VDPWR.n384 VDPWR.n370 5.78175
R3036 VDPWR.n259 VDPWR.n134 5.78175
R3037 VDPWR.n134 VDPWR.n105 5.78175
R3038 VDPWR.n264 VDPWR.n258 5.78175
R3039 VDPWR.n258 VDPWR.n113 5.78175
R3040 VDPWR.n257 VDPWR.n129 5.78175
R3041 VDPWR.n257 VDPWR.n113 5.78175
R3042 VDPWR.n290 VDPWR.n289 5.78175
R3043 VDPWR.n289 VDPWR.n105 5.78175
R3044 VDPWR.n130 VDPWR.n124 5.78175
R3045 VDPWR.n124 VDPWR.n115 5.78175
R3046 VDPWR.n297 VDPWR.n123 5.78175
R3047 VDPWR.n123 VDPWR.n115 5.78175
R3048 VDPWR.n206 VDPWR.n205 5.78175
R3049 VDPWR.n214 VDPWR.n206 5.78175
R3050 VDPWR.n216 VDPWR.n215 5.78175
R3051 VDPWR.n215 VDPWR.n214 5.78175
R3052 VDPWR.n121 VDPWR.n109 5.78175
R3053 VDPWR.n121 VDPWR.n115 5.78175
R3054 VDPWR.n140 VDPWR.n120 5.78175
R3055 VDPWR.n120 VDPWR.n115 5.78175
R3056 VDPWR.n191 VDPWR.n163 5.78175
R3057 VDPWR.n243 VDPWR.n163 5.78175
R3058 VDPWR.n192 VDPWR.n155 5.78175
R3059 VDPWR.n249 VDPWR.n155 5.78175
R3060 VDPWR.n248 VDPWR.n247 5.78175
R3061 VDPWR.n249 VDPWR.n248 5.78175
R3062 VDPWR.n245 VDPWR.n244 5.78175
R3063 VDPWR.n244 VDPWR.n243 5.78175
R3064 VDPWR.n279 VDPWR.n139 5.78175
R3065 VDPWR.n139 VDPWR.n105 5.78175
R3066 VDPWR.n269 VDPWR.n117 5.78175
R3067 VDPWR.n269 VDPWR.n113 5.78175
R3068 VDPWR.n274 VDPWR.n273 5.78175
R3069 VDPWR.n273 VDPWR.n113 5.78175
R3070 VDPWR.n276 VDPWR.n138 5.78175
R3071 VDPWR.n138 VDPWR.n105 5.78175
R3072 VDPWR.n239 VDPWR.n146 5.78175
R3073 VDPWR.n243 VDPWR.n146 5.78175
R3074 VDPWR.n235 VDPWR.n154 5.78175
R3075 VDPWR.n249 VDPWR.n154 5.78175
R3076 VDPWR.n236 VDPWR.n166 5.78175
R3077 VDPWR.n214 VDPWR.n166 5.78175
R3078 VDPWR.n253 VDPWR.n147 5.78175
R3079 VDPWR.n243 VDPWR.n147 5.78175
R3080 VDPWR.n251 VDPWR.n250 5.78175
R3081 VDPWR.n250 VDPWR.n249 5.78175
R3082 VDPWR.n170 VDPWR.n165 5.78175
R3083 VDPWR.n214 VDPWR.n165 5.78175
R3084 VDPWR.n583 VDPWR.n572 4.7119
R3085 VDPWR.n376 VDPWR.n362 4.7119
R3086 VDPWR.n342 VDPWR.n331 4.7119
R3087 VDPWR.n189 VDPWR.n185 4.7119
R3088 VDPWR.n228 VDPWR.n148 4.7119
R3089 VDPWR.n284 VDPWR.n278 4.7119
R3090 VDPWR.n135 VDPWR.n99 4.7119
R3091 VDPWR.n615 VDPWR.n614 4.70083
R3092 VDPWR.n387 VDPWR.n374 4.70083
R3093 VDPWR.n442 VDPWR.n441 4.70083
R3094 VDPWR.n199 VDPWR.n197 4.70083
R3095 VDPWR.n177 VDPWR.n176 4.70083
R3096 VDPWR.n119 VDPWR.n118 4.70083
R3097 VDPWR.n128 VDPWR.n127 4.70083
R3098 VDPWR.n625 VDPWR.n578 3.98297
R3099 VDPWR.n402 VDPWR.n401 3.98297
R3100 VDPWR.n452 VDPWR.n337 3.98297
R3101 VDPWR.n214 VDPWR.n213 3.98297
R3102 VDPWR.n115 VDPWR.n102 3.98297
R3103 VDPWR.n639 VDPWR 3.64817
R3104 VDPWR.n322 VDPWR 3.52106
R3105 VDPWR.n92 VDPWR 3.52106
R3106 VDPWR.n646 VDPWR.n645 3.32168
R3107 VDPWR VDPWR.n0 3.05185
R3108 VDPWR.n563 VDPWR 2.62366
R3109 VDPWR.n748 VDPWR 2.3405
R3110 VDPWR.n748 VDPWR 2.3405
R3111 VDPWR.n794 VDPWR 2.3405
R3112 VDPWR.n794 VDPWR 2.3405
R3113 VDPWR.n696 VDPWR 2.3405
R3114 VDPWR.n696 VDPWR 2.3405
R3115 VDPWR.n668 VDPWR 2.3405
R3116 VDPWR.n668 VDPWR 2.3405
R3117 VDPWR.n470 VDPWR 2.3405
R3118 VDPWR.n470 VDPWR 2.3405
R3119 VDPWR.n500 VDPWR 2.3405
R3120 VDPWR.n500 VDPWR 2.3405
R3121 VDPWR.n518 VDPWR 2.3405
R3122 VDPWR.n518 VDPWR 2.3405
R3123 VDPWR.n548 VDPWR 2.3405
R3124 VDPWR.n548 VDPWR 2.3405
R3125 VDPWR.n89 VDPWR 2.3405
R3126 VDPWR.n62 VDPWR 2.3405
R3127 VDPWR.n36 VDPWR 2.3405
R3128 VDPWR.n38 VDPWR 2.3405
R3129 VDPWR.n795 VDPWR 2.29412
R3130 VDPWR.n653 VDPWR 2.29412
R3131 VDPWR.n653 VDPWR 2.29412
R3132 VDPWR.n64 VDPWR 2.29412
R3133 VDPWR.n243 VDPWR.n242 1.99173
R3134 VDPWR.n281 VDPWR.n105 1.99173
R3135 VDPWR.n97 VDPWR 1.93224
R3136 VDPWR.n183 VDPWR 1.93224
R3137 VDPWR.n39 VDPWR.n38 1.92169
R3138 VDPWR.n459 VDPWR 1.89811
R3139 VDPWR.n407 VDPWR 1.89811
R3140 VDPWR.n749 VDPWR.n743 1.8605
R3141 VDPWR.n793 VDPWR.n731 1.8605
R3142 VDPWR.n697 VDPWR.n666 1.8605
R3143 VDPWR.n695 VDPWR.n667 1.8605
R3144 VDPWR.n750 VDPWR.n749 1.8605
R3145 VDPWR.n793 VDPWR.n792 1.8605
R3146 VDPWR.n698 VDPWR.n697 1.8605
R3147 VDPWR.n695 VDPWR.n694 1.8605
R3148 VDPWR.n510 VDPWR.n469 1.8605
R3149 VDPWR.n501 VDPWR.n499 1.8605
R3150 VDPWR.n510 VDPWR.n509 1.8605
R3151 VDPWR.n502 VDPWR.n501 1.8605
R3152 VDPWR.n558 VDPWR.n517 1.8605
R3153 VDPWR.n549 VDPWR.n547 1.8605
R3154 VDPWR.n558 VDPWR.n557 1.8605
R3155 VDPWR.n550 VDPWR.n549 1.8605
R3156 VDPWR.n37 VDPWR.n31 1.8605
R3157 VDPWR.n63 VDPWR.n11 1.8605
R3158 VDPWR.n88 VDPWR.n87 1.8605
R3159 VDPWR.n612 VDPWR.n610 1.77828
R3160 VDPWR.n439 VDPWR.n431 1.77828
R3161 VDPWR.n394 VDPWR.n393 1.77828
R3162 VDPWR.n194 VDPWR.n192 1.77828
R3163 VDPWR.n305 VDPWR.n117 1.77828
R3164 VDPWR.n299 VDPWR.n129 1.77828
R3165 VDPWR.n235 VDPWR.n234 1.77828
R3166 VDPWR.n834 VDPWR.n833 1.76063
R3167 VDPWR.n560 VDPWR.n559 1.76063
R3168 VDPWR.n464 VDPWR.n324 1.753
R3169 VDPWR.n644 VDPWR.n643 1.753
R3170 VDPWR.n512 VDPWR.n511 1.75125
R3171 VDPWR.n326 VDPWR.n325 1.603
R3172 VDPWR.n462 VDPWR.n461 1.603
R3173 VDPWR.n631 VDPWR 1.43984
R3174 VDPWR.n598 VDPWR.n596 1.3042
R3175 VDPWR.n353 VDPWR.n345 1.3042
R3176 VDPWR.n396 VDPWR.n395 1.3042
R3177 VDPWR.n217 VDPWR.n216 1.3042
R3178 VDPWR.n141 VDPWR.n140 1.3042
R3179 VDPWR.n131 VDPWR.n130 1.3042
R3180 VDPWR.n237 VDPWR.n236 1.3042
R3181 VDPWR.n589 VDPWR.n586 1.19372
R3182 VDPWR.n437 VDPWR.n436 1.19372
R3183 VDPWR.n391 VDPWR.n390 1.19372
R3184 VDPWR.n205 VDPWR.n188 1.19372
R3185 VDPWR.n313 VDPWR.n109 1.19372
R3186 VDPWR.n297 VDPWR.n296 1.19372
R3187 VDPWR.n174 VDPWR.n170 1.19372
R3188 VDPWR.n640 VDPWR.n3 1.18677
R3189 VDPWR.n833 VDPWR.n651 1.12394
R3190 VDPWR.n569 VDPWR.n465 1.10237
R3191 VDPWR.n511 VDPWR.n2 1.06531
R3192 VDPWR.n570 VDPWR 1.06379
R3193 VDPWR.n511 VDPWR.n510 1.06168
R3194 VDPWR.n559 VDPWR.n558 1.06168
R3195 VDPWR.n559 VDPWR.n516 1.05594
R3196 VDPWR.n329 VDPWR 1.04172
R3197 VDPWR.n411 VDPWR 1.04172
R3198 VDPWR.n321 VDPWR 0.890303
R3199 VDPWR.n182 VDPWR 0.890303
R3200 VDPWR.n568 VDPWR 0.859781
R3201 VDPWR.n458 VDPWR 0.854351
R3202 VDPWR.n406 VDPWR 0.854351
R3203 VDPWR.n562 VDPWR.n468 0.770146
R3204 VDPWR.n634 VDPWR 0.768852
R3205 VDPWR.n567 VDPWR 0.758767
R3206 VDPWR.n636 VDPWR.n635 0.73918
R3207 VDPWR.n831 VDPWR.n652 0.715885
R3208 VDPWR.n797 VDPWR.n796 0.715885
R3209 VDPWR.n831 VDPWR.n830 0.715885
R3210 VDPWR.n66 VDPWR.n65 0.715885
R3211 VDPWR.n408 VDPWR 0.69425
R3212 VDPWR.n460 VDPWR 0.69425
R3213 VDPWR.n562 VDPWR.n561 0.623777
R3214 VDPWR.n632 VDPWR.n631 0.619997
R3215 VDPWR.n570 VDPWR.n563 0.619997
R3216 VDPWR.n648 VDPWR.n90 0.615521
R3217 VDPWR.n90 VDPWR 0.559955
R3218 VDPWR.n97 VDPWR.n96 0.518921
R3219 VDPWR.n322 VDPWR.n321 0.518921
R3220 VDPWR.n183 VDPWR.n93 0.518921
R3221 VDPWR.n182 VDPWR.n92 0.518921
R3222 VDPWR.n639 VDPWR.n638 0.507812
R3223 VDPWR.n641 VDPWR.n640 0.507416
R3224 VDPWR.n95 VDPWR 0.505434
R3225 VDPWR.n645 VDPWR 0.505434
R3226 VDPWR.n329 VDPWR.n328 0.497975
R3227 VDPWR.n459 VDPWR.n458 0.497975
R3228 VDPWR.n407 VDPWR.n406 0.497975
R3229 VDPWR.n411 VDPWR.n410 0.497975
R3230 VDPWR.n646 VDPWR 0.467672
R3231 VDPWR.n323 VDPWR 0.467461
R3232 VDPWR VDPWR.n0 0.464224
R3233 VDPWR.n647 VDPWR.n646 0.426664
R3234 VDPWR.n796 VDPWR 0.413
R3235 VDPWR.n832 VDPWR.n831 0.410656
R3236 VDPWR.n694 VDPWR.n669 0.376971
R3237 VDPWR.n699 VDPWR.n698 0.376971
R3238 VDPWR.n830 VDPWR.n654 0.376971
R3239 VDPWR.n797 VDPWR.n730 0.376971
R3240 VDPWR.n792 VDPWR.n732 0.376971
R3241 VDPWR.n751 VDPWR.n750 0.376971
R3242 VDPWR.n675 VDPWR.n667 0.376971
R3243 VDPWR.n678 VDPWR.n666 0.376971
R3244 VDPWR.n820 VDPWR.n652 0.376971
R3245 VDPWR.n738 VDPWR.n731 0.376971
R3246 VDPWR.n744 VDPWR.n743 0.376971
R3247 VDPWR.n503 VDPWR.n502 0.376971
R3248 VDPWR.n509 VDPWR.n471 0.376971
R3249 VDPWR.n499 VDPWR.n482 0.376971
R3250 VDPWR.n492 VDPWR.n469 0.376971
R3251 VDPWR.n551 VDPWR.n550 0.376971
R3252 VDPWR.n557 VDPWR.n519 0.376971
R3253 VDPWR.n547 VDPWR.n530 0.376971
R3254 VDPWR.n540 VDPWR.n517 0.376971
R3255 VDPWR.n629 VDPWR.n571 0.376971
R3256 VDPWR.n456 VDPWR.n330 0.376971
R3257 VDPWR.n414 VDPWR.n413 0.376971
R3258 VDPWR.n87 VDPWR.n4 0.376971
R3259 VDPWR.n12 VDPWR.n11 0.376971
R3260 VDPWR.n67 VDPWR.n66 0.376971
R3261 VDPWR.n32 VDPWR.n31 0.376971
R3262 VDPWR.n40 VDPWR.n39 0.376971
R3263 VDPWR.n224 VDPWR.n184 0.376971
R3264 VDPWR.n110 VDPWR.n94 0.376971
R3265 VDPWR.n319 VDPWR.n98 0.376971
R3266 VDPWR.n226 VDPWR.n181 0.376971
R3267 VDPWR.n633 VDPWR 0.376726
R3268 VDPWR.n796 VDPWR.n795 0.360656
R3269 VDPWR.n831 VDPWR.n653 0.360656
R3270 VDPWR.n566 VDPWR 0.351319
R3271 VDPWR VDPWR.n568 0.345458
R3272 VDPWR.n635 VDPWR.n562 0.34097
R3273 VDPWR.n567 VDPWR.n566 0.327725
R3274 VDPWR.n566 VDPWR.n565 0.327725
R3275 VDPWR.n640 VDPWR.n639 0.321157
R3276 VDPWR.n613 VDPWR.n612 0.307571
R3277 VDPWR.n440 VDPWR.n439 0.307571
R3278 VDPWR.n393 VDPWR.n389 0.307571
R3279 VDPWR.n196 VDPWR.n194 0.307571
R3280 VDPWR.n305 VDPWR.n304 0.307571
R3281 VDPWR.n300 VDPWR.n299 0.307571
R3282 VDPWR.n234 VDPWR.n169 0.307571
R3283 VDPWR.n632 VDPWR 0.304352
R3284 VDPWR.n409 VDPWR 0.27355
R3285 VDPWR.n327 VDPWR 0.272663
R3286 VDPWR.n96 VDPWR 0.254776
R3287 VDPWR.n93 VDPWR 0.254776
R3288 VDPWR.n513 VDPWR.n512 0.249058
R3289 VDPWR.n463 VDPWR.n462 0.244984
R3290 VDPWR.n328 VDPWR 0.244503
R3291 VDPWR.n410 VDPWR 0.244503
R3292 VDPWR.n464 VDPWR.n463 0.234803
R3293 VDPWR.n561 VDPWR.n560 0.232427
R3294 VDPWR.n65 VDPWR.n0 0.22821
R3295 VDPWR.n515 VDPWR.n2 0.218931
R3296 VDPWR.n516 VDPWR.n468 0.204432
R3297 VDPWR.n65 VDPWR.n64 0.201986
R3298 VDPWR.n642 VDPWR.n465 0.193242
R3299 VDPWR.n512 VDPWR.n1 0.189404
R3300 VDPWR.n623 VDPWR.n622 0.178728
R3301 VDPWR.n450 VDPWR.n449 0.178728
R3302 VDPWR.n399 VDPWR.n398 0.178728
R3303 VDPWR.n191 VDPWR.n190 0.178728
R3304 VDPWR.n283 VDPWR.n279 0.178728
R3305 VDPWR.n290 VDPWR.n132 0.178728
R3306 VDPWR.n240 VDPWR.n239 0.178728
R3307 VDPWR.n651 VDPWR.n650 0.171208
R3308 VDPWR.n649 VDPWR.n3 0.171141
R3309 VDPWR.n648 VDPWR.n647 0.166741
R3310 VDPWR.n651 VDPWR.n2 0.166514
R3311 VDPWR.n697 VDPWR 0.166125
R3312 VDPWR.n793 VDPWR 0.164562
R3313 VDPWR VDPWR.n695 0.164562
R3314 VDPWR.n501 VDPWR 0.164562
R3315 VDPWR.n549 VDPWR 0.164562
R3316 VDPWR.n515 VDPWR.n514 0.163619
R3317 VDPWR.n468 VDPWR.n467 0.162949
R3318 VDPWR.n638 VDPWR.n637 0.153104
R3319 VDPWR.n641 VDPWR.n466 0.1514
R3320 VDPWR VDPWR.n460 0.148
R3321 VDPWR.n321 VDPWR.n320 0.147704
R3322 VDPWR.n225 VDPWR.n182 0.147704
R3323 VDPWR.n320 VDPWR.n97 0.146059
R3324 VDPWR.n225 VDPWR.n183 0.146059
R3325 VDPWR.n457 VDPWR.n456 0.133357
R3326 VDPWR.n413 VDPWR.n412 0.133357
R3327 VDPWR.n320 VDPWR.n94 0.133357
R3328 VDPWR.n320 VDPWR.n319 0.133357
R3329 VDPWR.n226 VDPWR.n225 0.133357
R3330 VDPWR.n225 VDPWR.n224 0.133357
R3331 VDPWR.n630 VDPWR.n629 0.133357
R3332 VDPWR.n96 VDPWR.n95 0.131257
R3333 VDPWR.n646 VDPWR.n92 0.131257
R3334 VDPWR.n645 VDPWR.n93 0.131257
R3335 VDPWR.n323 VDPWR.n322 0.129612
R3336 VDPWR.n636 VDPWR.n91 0.125788
R3337 VDPWR.n630 VDPWR.n570 0.110181
R3338 VDPWR.n749 VDPWR.n748 0.109875
R3339 VDPWR.n794 VDPWR.n793 0.109875
R3340 VDPWR.n697 VDPWR.n696 0.109875
R3341 VDPWR.n695 VDPWR.n668 0.109875
R3342 VDPWR.n510 VDPWR.n470 0.109875
R3343 VDPWR.n501 VDPWR.n500 0.109875
R3344 VDPWR.n558 VDPWR.n518 0.109875
R3345 VDPWR.n549 VDPWR.n548 0.109875
R3346 VDPWR.n564 VDPWR 0.109033
R3347 VDPWR.n631 VDPWR.n630 0.108956
R3348 VDPWR VDPWR.n323 0.100037
R3349 VDPWR.n633 VDPWR.n632 0.0979265
R3350 VDPWR.n623 VDPWR.n582 0.0977152
R3351 VDPWR.n450 VDPWR.n341 0.0977152
R3352 VDPWR.n398 VDPWR.n397 0.0977152
R3353 VDPWR.n218 VDPWR.n191 0.0977152
R3354 VDPWR.n279 VDPWR.n108 0.0977152
R3355 VDPWR.n291 VDPWR.n290 0.0977152
R3356 VDPWR.n239 VDPWR.n238 0.0977152
R3357 VDPWR.n634 VDPWR.n563 0.096701
R3358 VDPWR.n564 VDPWR 0.0963995
R3359 VDPWR.n565 VDPWR 0.096377
R3360 VDPWR.n514 VDPWR.n513 0.0952222
R3361 VDPWR.n650 VDPWR.n1 0.0952222
R3362 VDPWR.n561 VDPWR.n467 0.0952222
R3363 VDPWR VDPWR.n63 0.0931573
R3364 VDPWR VDPWR.n37 0.0922832
R3365 VDPWR.n88 VDPWR 0.0922832
R3366 VDPWR.n650 VDPWR.n649 0.0884817
R3367 VDPWR.n458 VDPWR.n457 0.079844
R3368 VDPWR.n412 VDPWR.n406 0.079844
R3369 VDPWR.n514 VDPWR.n466 0.0789784
R3370 VDPWR.n457 VDPWR.n329 0.0789574
R3371 VDPWR.n412 VDPWR.n411 0.0789574
R3372 VDPWR.n637 VDPWR.n467 0.078882
R3373 VDPWR.n833 VDPWR.n832 0.0780862
R3374 VDPWR.n834 VDPWR.n1 0.0742538
R3375 VDPWR.n638 VDPWR.n465 0.0715417
R3376 VDPWR.n328 VDPWR.n327 0.0709787
R3377 VDPWR.n460 VDPWR.n459 0.0709787
R3378 VDPWR.n408 VDPWR.n407 0.0709787
R3379 VDPWR.n410 VDPWR.n409 0.0700922
R3380 VDPWR.n569 VDPWR 0.0630773
R3381 VDPWR.n643 VDPWR.n642 0.0627018
R3382 VDPWR.n463 VDPWR.n3 0.0625
R3383 VDPWR.n37 VDPWR.n36 0.0616888
R3384 VDPWR.n63 VDPWR.n62 0.0616888
R3385 VDPWR.n89 VDPWR.n88 0.0616888
R3386 VDPWR.n642 VDPWR.n641 0.0573333
R3387 VDPWR.n635 VDPWR.n634 0.0572867
R3388 VDPWR.n748 VDPWR 0.0551875
R3389 VDPWR VDPWR.n794 0.0551875
R3390 VDPWR.n696 VDPWR 0.0551875
R3391 VDPWR.n668 VDPWR 0.0551875
R3392 VDPWR VDPWR.n470 0.0551875
R3393 VDPWR.n500 VDPWR 0.0551875
R3394 VDPWR VDPWR.n518 0.0551875
R3395 VDPWR.n548 VDPWR 0.0551875
R3396 VDPWR.n647 VDPWR.n91 0.0549669
R3397 VDPWR.n461 VDPWR 0.0545625
R3398 VDPWR.n795 VDPWR 0.0512812
R3399 VDPWR VDPWR.n653 0.0512812
R3400 VDPWR.n633 VDPWR.n569 0.045162
R3401 VDPWR.n649 VDPWR.n648 0.043125
R3402 VDPWR.n637 VDPWR.n636 0.03925
R3403 VDPWR.n643 VDPWR.n464 0.0388531
R3404 VDPWR.n466 VDPWR.n91 0.0360208
R3405 VDPWR.n409 VDPWR.n326 0.0351875
R3406 VDPWR.n324 VDPWR 0.0334335
R3407 VDPWR.n645 VDPWR.n644 0.0315396
R3408 VDPWR.n38 VDPWR 0.0310944
R3409 VDPWR.n36 VDPWR 0.0310944
R3410 VDPWR.n62 VDPWR 0.0310944
R3411 VDPWR VDPWR.n89 0.0310944
R3412 VDPWR.n408 VDPWR.n90 0.0298951
R3413 VDPWR.n64 VDPWR 0.0289091
R3414 VDPWR.n327 VDPWR 0.0265417
R3415 VDPWR.n462 VDPWR.n325 0.0256039
R3416 VDPWR.n560 VDPWR.n513 0.0160462
R3417 VDPWR.n516 VDPWR.n515 0.0149983
R3418 VDPWR.n95 VDPWR 0.0140031
R3419 VDPWR.n461 VDPWR.n326 0.008
R3420 VDPWR.n95 VDPWR 0.00744444
R3421 VDPWR VDPWR.n834 0.00538077
R3422 VDPWR.n325 VDPWR 0.00308012
R3423 VDPWR.n832 VDPWR 0.00284375
R3424 VDPWR.n565 VDPWR.n564 0.00149206
R3425 VDPWR.n568 VDPWR.n567 0.00149206
R3426 VDPWR.n644 VDPWR.n324 0.00113131
R3427 ua[1].n1 ua[1] 9.55241
R3428 ua[1].n0 ua[1] 2.51601
R3429 ua[1].n0 ua[1] 2.11902
R3430 ua[1].n1 ua[1].n0 0.188289
R3431 ua[1] ua[1].n1 0.0879542
R3432 flashADC_3bit_0/comp_p_1/out_left.n1 flashADC_3bit_0/comp_p_1/out_left.t2 145.612
R3433 flashADC_3bit_0/comp_p_1/out_left.n2 flashADC_3bit_0/comp_p_1/out_left.t0 143.417
R3434 flashADC_3bit_0/comp_p_1/out_left.n0 flashADC_3bit_0/comp_p_1/out_left.t1 29.4286
R3435 flashADC_3bit_0/comp_p_1/out_left flashADC_3bit_0/comp_p_1/out_left.n3 11.6041
R3436 flashADC_3bit_0/comp_p_1/out_left.n3 flashADC_3bit_0/comp_p_1/out_left.n2 4.33076
R3437 flashADC_3bit_0/comp_p_1/out_left.n1 flashADC_3bit_0/comp_p_1/out_left.n0 2.12634
R3438 flashADC_3bit_0/comp_p_1/out_left.n2 flashADC_3bit_0/comp_p_1/out_left.n1 2.04428
R3439 flashADC_3bit_0/comp_p_1/out_left.n3 flashADC_3bit_0/comp_p_1/out_left.n0 0.00290385
R3440 uo_out[3].n0 uo_out[3].t1 556.78
R3441 uo_out[3].t1 uo_out[3] 547.24
R3442 uo_out[3] uo_out[3].t0 372.113
R3443 uo_out[3].n0 uo_out[3] 9.54008
R3444 uo_out[3].n3 uo_out[3].n2 4.55415
R3445 uo_out[3].n2 uo_out[3] 4.43618
R3446 uo_out[3].n3 uo_out[3] 3.33965
R3447 uo_out[3].n1 uo_out[3].n0 0.253625
R3448 uo_out[3] uo_out[3] 0.063
R3449 uo_out[3].n2 uo_out[3] 0.0443144
R3450 uo_out[3] uo_out[3].n3 0.0262742
R3451 uo_out[3] uo_out[3] 0.0262732
R3452 uo_out[3].n1 uo_out[3] 0.013
R3453 uo_out[3].n3 uo_out[3] 0.00801031
R3454 uo_out[3] uo_out[3].n1 0.00565464
R3455 ua[0].n20 ua[0].t26 899.324
R3456 ua[0].n38 ua[0].t22 899.324
R3457 ua[0].n31 ua[0].t14 899.324
R3458 ua[0].n25 ua[0].t2 899.324
R3459 ua[0].n2 ua[0].t6 899.324
R3460 ua[0].n7 ua[0].t10 899.324
R3461 ua[0].n13 ua[0].t18 899.324
R3462 ua[0].n21 ua[0].t26 898.659
R3463 ua[0].n39 ua[0].t22 898.659
R3464 ua[0].n32 ua[0].t14 898.659
R3465 ua[0].n26 ua[0].t2 898.659
R3466 ua[0].n3 ua[0].t6 898.659
R3467 ua[0].n8 ua[0].t10 898.659
R3468 ua[0].n14 ua[0].t18 898.659
R3469 ua[0].t23 ua[0].n38 898.442
R3470 ua[0].t3 ua[0].n25 898.442
R3471 ua[0].t7 ua[0].n2 898.442
R3472 ua[0].t19 ua[0].n13 898.442
R3473 ua[0].t27 ua[0].n20 898.442
R3474 ua[0].t15 ua[0].n31 898.442
R3475 ua[0].t11 ua[0].n7 898.442
R3476 ua[0].n21 ua[0].t27 897.754
R3477 ua[0].n39 ua[0].t23 897.754
R3478 ua[0].n32 ua[0].t15 897.754
R3479 ua[0].n26 ua[0].t3 897.754
R3480 ua[0].n3 ua[0].t7 897.754
R3481 ua[0].n8 ua[0].t11 897.754
R3482 ua[0].n14 ua[0].t19 897.754
R3483 ua[0].n18 ua[0].t24 895.625
R3484 ua[0].n36 ua[0].t20 895.625
R3485 ua[0].n29 ua[0].t12 895.625
R3486 ua[0].n23 ua[0].t0 895.625
R3487 ua[0].n0 ua[0].t4 895.625
R3488 ua[0].n5 ua[0].t8 895.625
R3489 ua[0].n11 ua[0].t16 895.625
R3490 ua[0].n18 ua[0].t25 894.172
R3491 ua[0].n36 ua[0].t21 894.172
R3492 ua[0].n29 ua[0].t13 894.172
R3493 ua[0].n23 ua[0].t1 894.172
R3494 ua[0].n0 ua[0].t5 894.172
R3495 ua[0].n5 ua[0].t9 894.172
R3496 ua[0].n11 ua[0].t17 894.172
R3497 ua[0] ua[0] 11.363
R3498 ua[0].n19 ua[0].n18 6.30807
R3499 ua[0].n37 ua[0].n36 6.30807
R3500 ua[0].n30 ua[0].n29 6.30807
R3501 ua[0].n24 ua[0].n23 6.30807
R3502 ua[0].n1 ua[0].n0 6.30807
R3503 ua[0].n6 ua[0].n5 6.30807
R3504 ua[0].n12 ua[0].n11 6.30807
R3505 ua[0].n20 ua[0].n19 5.39021
R3506 ua[0].n38 ua[0].n37 5.39021
R3507 ua[0].n31 ua[0].n30 5.39021
R3508 ua[0].n25 ua[0].n24 5.39021
R3509 ua[0].n2 ua[0].n1 5.39021
R3510 ua[0].n7 ua[0].n6 5.39021
R3511 ua[0].n13 ua[0].n12 5.39021
R3512 ua[0].n22 ua[0].n21 5.38653
R3513 ua[0].n40 ua[0].n39 5.38653
R3514 ua[0].n33 ua[0].n32 5.38653
R3515 ua[0].n27 ua[0].n26 5.38653
R3516 ua[0].n4 ua[0].n3 5.38653
R3517 ua[0].n9 ua[0].n8 5.38653
R3518 ua[0].n15 ua[0].n14 5.38653
R3519 ua[0].n44 ua[0].n43 5.20469
R3520 ua[0].n22 ua[0].n19 5.11108
R3521 ua[0].n40 ua[0].n37 5.11108
R3522 ua[0].n33 ua[0].n30 5.11108
R3523 ua[0].n27 ua[0].n24 5.11108
R3524 ua[0].n4 ua[0].n1 5.11108
R3525 ua[0].n9 ua[0].n6 5.11108
R3526 ua[0].n15 ua[0].n12 5.11108
R3527 ua[0].n35 ua[0].n28 4.57467
R3528 ua[0].n10 ua[0] 4.13219
R3529 ua[0].n35 ua[0].n34 3.68222
R3530 ua[0].n42 ua[0].n41 3.10272
R3531 ua[0].n16 ua[0] 2.68025
R3532 ua[0].n10 ua[0] 2.66582
R3533 ua[0].n43 ua[0].n42 2.43775
R3534 ua[0].n43 ua[0] 1.54614
R3535 ua[0].n17 ua[0].n16 1.35915
R3536 ua[0] ua[0].n22 0.870692
R3537 ua[0] ua[0].n4 0.870692
R3538 ua[0] ua[0].n9 0.870692
R3539 ua[0] ua[0].n15 0.870692
R3540 ua[0].n34 ua[0].n33 0.837038
R3541 ua[0].n41 ua[0].n40 0.726462
R3542 ua[0].n16 ua[0].n10 0.70492
R3543 ua[0].n28 ua[0].n27 0.668769
R3544 ua[0].n42 ua[0].n35 0.533734
R3545 ua[0].n17 ua[0] 0.468179
R3546 ua[0] ua[0].n45 0.332981
R3547 ua[0].n45 ua[0] 0.20608
R3548 ua[0].n41 ua[0] 0.0482941
R3549 ua[0].n44 ua[0].n17 0.0422977
R3550 ua[0].n45 ua[0].n44 0.0422977
R3551 ua[0].n28 ua[0] 0.0391905
R3552 ua[0].n34 ua[0] 0.0341538
R3553 flashADC_3bit_0/comp_p_0/latch_left.n0 flashADC_3bit_0/comp_p_0/latch_left.t3 114.778
R3554 flashADC_3bit_0/comp_p_0/latch_left.n0 flashADC_3bit_0/comp_p_0/latch_left.t2 106.572
R3555 flashADC_3bit_0/comp_p_0/latch_left.n1 flashADC_3bit_0/comp_p_0/latch_left.t0 95.1712
R3556 flashADC_3bit_0/comp_p_0/latch_left.n2 flashADC_3bit_0/comp_p_0/latch_left.t1 22.0141
R3557 flashADC_3bit_0/comp_p_0/latch_left.n1 flashADC_3bit_0/comp_p_0/latch_left.n0 1.72733
R3558 flashADC_3bit_0/comp_p_0/latch_left flashADC_3bit_0/comp_p_0/latch_left.n2 0.717514
R3559 flashADC_3bit_0/comp_p_0/latch_left.n2 flashADC_3bit_0/comp_p_0/latch_left.n1 0.599169
R3560 uo_out[4].n0 uo_out[4].t1 556.78
R3561 uo_out[4].t1 uo_out[4] 547.24
R3562 uo_out[4] uo_out[4].t0 372.113
R3563 uo_out[4].n1 uo_out[4] 20.4931
R3564 uo_out[4].n0 uo_out[4] 9.54008
R3565 uo_out[4].n2 uo_out[4] 4.35598
R3566 uo_out[4].n2 uo_out[4].n1 3.45922
R3567 uo_out[4].n1 uo_out[4] 1.38807
R3568 uo_out[4] uo_out[4].n0 0.266125
R3569 uo_out[4] uo_out[4] 0.063
R3570 uo_out[4] uo_out[4].n2 0.0217258
R3571 uo_out[4].n2 uo_out[4] 0.00887356
R3572 flashADC_3bit_0/comp_p_2/out_left.n1 flashADC_3bit_0/comp_p_2/out_left.t2 145.612
R3573 flashADC_3bit_0/comp_p_2/out_left.n2 flashADC_3bit_0/comp_p_2/out_left.t0 143.417
R3574 flashADC_3bit_0/comp_p_2/out_left.n0 flashADC_3bit_0/comp_p_2/out_left.t1 29.4286
R3575 flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/comp_p_2/out_left.n3 11.6041
R3576 flashADC_3bit_0/comp_p_2/out_left.n3 flashADC_3bit_0/comp_p_2/out_left.n2 4.33076
R3577 flashADC_3bit_0/comp_p_2/out_left.n1 flashADC_3bit_0/comp_p_2/out_left.n0 2.12634
R3578 flashADC_3bit_0/comp_p_2/out_left.n2 flashADC_3bit_0/comp_p_2/out_left.n1 2.04428
R3579 flashADC_3bit_0/comp_p_2/out_left.n3 flashADC_3bit_0/comp_p_2/out_left.n0 0.00290385
R3580 uo_out[5].n0 uo_out[5].t1 556.78
R3581 uo_out[5].t1 uo_out[5] 547.24
R3582 uo_out[5] uo_out[5].t0 372.113
R3583 uo_out[5].n2 uo_out[5] 18.5756
R3584 uo_out[5].n0 uo_out[5] 9.54008
R3585 uo_out[5].n3 uo_out[5] 5.91776
R3586 uo_out[5].n2 uo_out[5] 1.06075
R3587 uo_out[5].n3 uo_out[5].n2 0.928508
R3588 uo_out[5].n1 uo_out[5].n0 0.25675
R3589 uo_out[5] uo_out[5].n3 0.0929839
R3590 uo_out[5] uo_out[5] 0.063
R3591 uo_out[5] uo_out[5] 0.0329675
R3592 uo_out[5].n3 uo_out[5] 0.0124426
R3593 uo_out[5].n1 uo_out[5] 0.009875
R3594 uo_out[5] uo_out[5].n1 0.00537013
R3595 flashADC_3bit_0/comp_p_3/latch_left.n0 flashADC_3bit_0/comp_p_3/latch_left.t3 114.778
R3596 flashADC_3bit_0/comp_p_3/latch_left.n0 flashADC_3bit_0/comp_p_3/latch_left.t2 106.572
R3597 flashADC_3bit_0/comp_p_3/latch_left.n1 flashADC_3bit_0/comp_p_3/latch_left.t0 95.1712
R3598 flashADC_3bit_0/comp_p_3/latch_left.n2 flashADC_3bit_0/comp_p_3/latch_left.t1 22.0141
R3599 flashADC_3bit_0/comp_p_3/latch_left.n1 flashADC_3bit_0/comp_p_3/latch_left.n0 1.72733
R3600 flashADC_3bit_0/comp_p_3/latch_left flashADC_3bit_0/comp_p_3/latch_left.n2 0.717514
R3601 flashADC_3bit_0/comp_p_3/latch_left.n2 flashADC_3bit_0/comp_p_3/latch_left.n1 0.599169
R3602 flashADC_3bit_0/comp_p_3/out_left.n1 flashADC_3bit_0/comp_p_3/out_left.t2 145.612
R3603 flashADC_3bit_0/comp_p_3/out_left.n2 flashADC_3bit_0/comp_p_3/out_left.t0 143.417
R3604 flashADC_3bit_0/comp_p_3/out_left.n0 flashADC_3bit_0/comp_p_3/out_left.t1 29.4286
R3605 flashADC_3bit_0/comp_p_3/out_left flashADC_3bit_0/comp_p_3/out_left.n3 11.6041
R3606 flashADC_3bit_0/comp_p_3/out_left.n3 flashADC_3bit_0/comp_p_3/out_left.n2 4.33076
R3607 flashADC_3bit_0/comp_p_3/out_left.n1 flashADC_3bit_0/comp_p_3/out_left.n0 2.12634
R3608 flashADC_3bit_0/comp_p_3/out_left.n2 flashADC_3bit_0/comp_p_3/out_left.n1 2.04428
R3609 flashADC_3bit_0/comp_p_3/out_left.n3 flashADC_3bit_0/comp_p_3/out_left.n0 0.00290385
R3610 uo_out[6].n0 uo_out[6].t1 556.78
R3611 uo_out[6].t1 uo_out[6] 547.24
R3612 uo_out[6] uo_out[6].t0 372.113
R3613 uo_out[6].n1 uo_out[6] 10.0074
R3614 uo_out[6].n0 uo_out[6] 9.54008
R3615 uo_out[6].n3 uo_out[6] 7.20627
R3616 uo_out[6].n2 uo_out[6].n1 1.978
R3617 uo_out[6].n1 uo_out[6] 0.589103
R3618 uo_out[6] uo_out[6].n0 0.266125
R3619 uo_out[6] uo_out[6].n3 0.0975323
R3620 uo_out[6] uo_out[6] 0.063
R3621 uo_out[6].n3 uo_out[6].n2 0.0223063
R3622 uo_out[6].n2 uo_out[6] 0.00579279
R3623 flashADC_3bit_0/comp_p_4/out_left.n1 flashADC_3bit_0/comp_p_4/out_left.t2 145.612
R3624 flashADC_3bit_0/comp_p_4/out_left.n2 flashADC_3bit_0/comp_p_4/out_left.t0 143.417
R3625 flashADC_3bit_0/comp_p_4/out_left.n0 flashADC_3bit_0/comp_p_4/out_left.t1 29.4286
R3626 flashADC_3bit_0/comp_p_4/out_left flashADC_3bit_0/comp_p_4/out_left.n3 11.6041
R3627 flashADC_3bit_0/comp_p_4/out_left.n3 flashADC_3bit_0/comp_p_4/out_left.n2 4.33076
R3628 flashADC_3bit_0/comp_p_4/out_left.n1 flashADC_3bit_0/comp_p_4/out_left.n0 2.12634
R3629 flashADC_3bit_0/comp_p_4/out_left.n2 flashADC_3bit_0/comp_p_4/out_left.n1 2.04428
R3630 flashADC_3bit_0/comp_p_4/out_left.n3 flashADC_3bit_0/comp_p_4/out_left.n0 0.00290385
R3631 uo_out[7].n0 uo_out[7].t1 556.78
R3632 uo_out[7].t1 uo_out[7] 547.24
R3633 uo_out[7] uo_out[7].t0 372.113
R3634 uo_out[7].n1 uo_out[7] 24.2927
R3635 uo_out[7].n0 uo_out[7] 9.54008
R3636 uo_out[7].n2 uo_out[7] 8.84384
R3637 uo_out[7].n1 uo_out[7] 1.81119
R3638 uo_out[7].n2 uo_out[7].n1 1.17633
R3639 uo_out[7] uo_out[7].n0 0.266125
R3640 uo_out[7] uo_out[7] 0.063
R3641 uo_out[7].n2 uo_out[7] 0.0115379
R3642 uo_out[7] uo_out[7].n2 0.00656452
R3643 uio_out[0].n0 uio_out[0].t1 556.78
R3644 uio_out[0].t1 uio_out[0] 547.24
R3645 uio_out[0] uio_out[0].t0 372.113
R3646 uio_out[0].n2 uio_out[0] 9.82897
R3647 uio_out[0].n0 uio_out[0] 9.54008
R3648 uio_out[0].n2 uio_out[0].n1 3.01518
R3649 uio_out[0].n1 uio_out[0] 2.80934
R3650 uio_out[0].n1 uio_out[0] 0.322375
R3651 uio_out[0] uio_out[0].n0 0.266125
R3652 uio_out[0] uio_out[0] 0.063
R3653 uio_out[0] uio_out[0].n2 0.0213143
R3654 flashADC_3bit_0/comp_p_6/out_left.n1 flashADC_3bit_0/comp_p_6/out_left.t2 145.612
R3655 flashADC_3bit_0/comp_p_6/out_left.n2 flashADC_3bit_0/comp_p_6/out_left.t0 143.417
R3656 flashADC_3bit_0/comp_p_6/out_left.n0 flashADC_3bit_0/comp_p_6/out_left.t1 29.4286
R3657 flashADC_3bit_0/comp_p_6/out_left flashADC_3bit_0/comp_p_6/out_left.n3 11.6041
R3658 flashADC_3bit_0/comp_p_6/out_left.n3 flashADC_3bit_0/comp_p_6/out_left.n2 4.33076
R3659 flashADC_3bit_0/comp_p_6/out_left.n1 flashADC_3bit_0/comp_p_6/out_left.n0 2.12634
R3660 flashADC_3bit_0/comp_p_6/out_left.n2 flashADC_3bit_0/comp_p_6/out_left.n1 2.04428
R3661 flashADC_3bit_0/comp_p_6/out_left.n3 flashADC_3bit_0/comp_p_6/out_left.n0 0.00290385
R3662 uio_out[1].n0 uio_out[1].t1 556.78
R3663 uio_out[1].t1 uio_out[1] 547.24
R3664 uio_out[1] uio_out[1].t0 372.113
R3665 uio_out[1].n1 uio_out[1] 11.4942
R3666 uio_out[1].n2 uio_out[1] 11.3634
R3667 uio_out[1].n0 uio_out[1] 9.54008
R3668 uio_out[1].n2 uio_out[1].n1 3.83483
R3669 uio_out[1].n1 uio_out[1] 1.33473
R3670 uio_out[1] uio_out[1].n0 0.266125
R3671 uio_out[1] uio_out[1] 0.063
R3672 uio_out[1] uio_out[1].n2 0.0550806
R3673 uio_out[1].n2 uio_out[1] 0.0207361
R3674 uo_out[0].n0 uo_out[0] 8.08738
R3675 uo_out[0].n0 uo_out[0] 5.30089
R3676 uo_out[0].n0 uo_out[0] 2.61734
R3677 uo_out[0] uo_out[0].n0 0.03175
R3678 uo_out[1].n0 uo_out[1] 9.67858
R3679 uo_out[1].n0 uo_out[1] 5.30089
R3680 uo_out[1].n0 uo_out[1] 2.61734
R3681 uo_out[1] uo_out[1].n0 0.03175
R3682 uo_out[2].n0 uo_out[2] 11.1559
R3683 uo_out[2].n0 uo_out[2] 5.30089
R3684 uo_out[2].n0 uo_out[2] 2.61734
R3685 uo_out[2] uo_out[2].n0 0.03175
C0 ua[6] ua[1] 0.01737f
C1 flashADC_3bit_0/comp_p_5/latch_left VDPWR 0.38506f
C2 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_4/vinn -0.04257f
C3 VDPWR flashADC_3bit_0/comp_p_5/out_left 0.47743f
C4 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_3/vinn -0.01472f
C5 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0.01085f
C6 uio_oe[3] uio_oe[4] 0.03102f
C7 ui_in[7] ui_in[6] 0.03102f
C8 uio_oe[2] VDPWR 0
C9 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G uo_out[2] 0
C10 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/m1_n100_n100# VDPWR 0.00545f
C11 uo_out[7] uio_out[1] 0
C12 uio_out[7] uio_out[6] 0.03102f
C13 uo_out[6] uo_out[7] 0.83703f
C14 ui_in[1] ui_in[2] 0.03102f
C15 flashADC_3bit_0/comp_p_5/vinn uo_out[7] -0.01219f
C16 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A 0.00574f
C17 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out uo_out[0] 0
C18 uo_out[5] uio_out[1] 0
C19 VDPWR uio_out[1] 2.03753f
C20 uo_out[6] uo_out[5] 0.83351f
C21 uo_out[6] VDPWR 0.59661f
C22 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 0.87869f
C23 uo_out[1] flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 0
C24 VDPWR flashADC_3bit_0/comp_p_2/tail 0.00107f
C25 flashADC_3bit_0/comp_p_3/latch_right VDPWR 0.26506f
C26 flashADC_3bit_0/comp_p_5/vinn VDPWR 3.18346f
C27 VDPWR flashADC_3bit_0/comp_p_0/out_left 0.12984f
C28 uio_out[2] VDPWR 0
C29 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_0/vinn -0.00292f
C30 ua[5] ua[1] 0.01737f
C31 uo_out[3] uo_out[0] 0
C32 VDPWR flashADC_3bit_0/comp_p_3/latch_left 0.27789f
C33 flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_0/vinn -0.03853f
C34 uio_in[3] uo_out[2] 0.00766f
C35 uio_oe[1] VDPWR 0
C36 VDPWR flashADC_3bit_0/comp_p_2/latch_right 0.23507f
C37 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A uo_out[2] 0
C38 uo_out[6] uo_out[2] 0
C39 uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 0.00393f
C40 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G VDPWR 0.10354f
C41 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G VDPWR 0.01001f
C42 uio_in[7] VDPWR 0
C43 ua[1] VDPWR 0.29111f
C44 VDPWR flashADC_3bit_0/comp_p_6/vinn 0.75805f
C45 flashADC_3bit_0/comp_p_4/latch_left VDPWR 0.25376f
C46 VDPWR flashADC_3bit_0/comp_p_4/tail 0.66705f
C47 flashADC_3bit_0/comp_p_0/tail VDPWR 0
C48 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin uo_out[1] 0.00143f
C49 uio_oe[0] VDPWR 0
C50 uo_out[4] uo_out[3] 0.31058f
C51 flashADC_3bit_0/comp_p_4/vinn ua[0] -0
C52 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_0/out_left -0.00559f
C53 uio_out[0] uio_out[1] 0.94888f
C54 uo_out[6] uio_out[0] 0
C55 flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_2/tail -0.01138f
C56 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_3/vinn -0.02012f
C57 uio_out[6] uio_out[5] 0.03102f
C58 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B -0
C59 uio_oe[3] uio_oe[2] 0.03102f
C60 ui_in[5] ui_in[6] 0.03102f
C61 uo_out[7] ua[0] -0
C62 uio_in[4] uio_in[3] 0.03102f
C63 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_2/latch_right -0.00771f
C64 uio_in[6] VDPWR 0
C65 ui_in[1] ui_in[0] 0.03102f
C66 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin uo_out[2] 0
C67 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin uo_out[5] 0
C68 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin VDPWR 0.01579f
C69 flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_2/latch_right -0.01316f
C70 VDPWR flashADC_3bit_0/comp_p_6/tail 0.00165f
C71 VDPWR ua[0] 6.62902f
C72 uio_in[6] uio_in[5] 0.03102f
C73 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin VDPWR 0.0018f
C74 flashADC_3bit_0/comp_p_1/tail VDPWR 0.02796f
C75 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 VDPWR 0.0044f
C76 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in 0
C77 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in 0.01474f
C78 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in uo_out[1] 0.00251f
C79 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin VDPWR 0.0016f
C80 VDPWR flashADC_3bit_0/comp_p_5/tail 0.78378f
C81 uio_out[7] VDPWR 0
C82 VDPWR flashADC_3bit_0/comp_p_3/tail 0.03261f
C83 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out VDPWR 1.04758f
C84 uio_out[3] uio_out[2] 0.03102f
C85 uo_out[0] uo_out[1] 1.70165f
C86 VDPWR uo_out[0] 0.10165f
C87 VDPWR flashADC_3bit_0/comp_p_4/latch_right 0.29499f
C88 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out 0.12659f
C89 VDPWR flashADC_3bit_0/comp_p_0/latch_left 0.16971f
C90 flashADC_3bit_0/comp_p_6/latch_left VDPWR 0.42219f
C91 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in uo_out[2] 0
C92 uio_in[5] uo_out[0] 0.01741f
C93 VDPWR flashADC_3bit_0/comp_p_5/latch_right 0.3836f
C94 uio_out[5] uio_out[4] 0.03102f
C95 flashADC_3bit_0/comp_p_1/latch_left VDPWR 0.23151f
C96 uo_out[6] uio_out[1] 0
C97 flashADC_3bit_0/comp_p_1/vinn ua[0] -0.00683f
C98 uio_oe[2] uio_oe[1] 0.03102f
C99 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out VDPWR 0.45869f
C100 uo_out[0] uo_out[2] 0.0867f
C101 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out uo_out[1] 0
C102 flashADC_3bit_0/comp_p_0/latch_right VDPWR 0.19561f
C103 uio_out[6] VDPWR 0
C104 uo_out[3] uo_out[7] 0
C105 uio_out[2] uio_out[1] 0.03102f
C106 flashADC_3bit_0/comp_p_3/vinn ua[0] -0.02041f
C107 uio_oe[7] uio_oe[6] 0.03102f
C108 flashADC_3bit_0/comp_p_4/out_left VDPWR 0.36618f
C109 uio_in[3] uio_in[2] 0.03102f
C110 flashADC_3bit_0/comp_p_2/vinn VDPWR 0.04885f
C111 uo_out[4] uo_out[7] 0
C112 ui_in[0] rst_n 0.03102f
C113 ua[1] ua[4] 0.01737f
C114 uo_out[3] uo_out[1] 0
C115 uo_out[3] uo_out[5] 0
C116 uo_out[3] VDPWR 0.20792f
C117 flashADC_3bit_0/comp_p_2/latch_left VDPWR 0.20391f
C118 ui_in[5] ui_in[4] 0.03102f
C119 uo_out[4] VDPWR 0.65166f
C120 uo_out[4] uo_out[5] 0.69387f
C121 flashADC_3bit_0/comp_p_6/vbias_p VDPWR 5.47005f
C122 flashADC_3bit_0/comp_p_1/out_left uo_out[7] 0
C123 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out uo_out[2] 0
C124 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_0/latch_left -0.01177f
C125 flashADC_3bit_0/comp_p_0/vinn ua[0] -0
C126 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out 0.00956f
C127 flashADC_3bit_0/comp_p_1/out_left VDPWR 0.15235f
C128 uo_out[3] uo_out[2] 0.09111f
C129 uio_out[5] VDPWR 0
C130 uio_oe[7] VDPWR 0
C131 uo_out[4] uo_out[2] 0
C132 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_6/vinn -0.01917f
C133 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_4/latch_left -0.02278f
C134 ua[1] ua[3] 0.01737f
C135 uio_in[1] uio_in[2] 0.03102f
C136 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_4/tail -0.04111f
C137 flashADC_3bit_0/comp_p_0/latch_right flashADC_3bit_0/comp_p_1/vinn -0.0159f
C138 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin VDPWR 0.00218f
C139 flashADC_3bit_0/comp_p_2/latch_left flashADC_3bit_0/comp_p_1/vinn -0.00559f
C140 flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_3/vinn -0.01451f
C141 uio_out[0] uo_out[3] 0.00111f
C142 uio_oe[1] uio_oe[0] 0.03102f
C143 uio_out[4] VDPWR 0
C144 flashADC_3bit_0/comp_p_2/latch_left flashADC_3bit_0/comp_p_3/vinn -0.00981f
C145 uo_out[4] flashADC_3bit_0/comp_p_1/vinn -0.01018f
C146 flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_1/vinn -0.00683f
C147 uio_oe[6] uio_oe[5] 0.03102f
C148 uio_oe[6] VDPWR 0
C149 uo_out[4] flashADC_3bit_0/comp_p_3/vinn -0
C150 flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_3/vinn -0.02616f
C151 flashADC_3bit_0/comp_p_6/vbias_p uio_out[0] 0
C152 rst_n clk 0.03102f
C153 ua[1] ua[2] 0.01737f
C154 flashADC_3bit_0/comp_p_5/vinn ua[0] -0.04026f
C155 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B 0.21063f
C156 uo_out[1] flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B 0
C157 flashADC_3bit_0/comp_p_1/tail uio_out[1] 0
C158 ui_in[4] ui_in[3] 0.03102f
C159 flashADC_3bit_0/comp_p_4/vinn VDPWR 0.57174f
C160 ua[1] flashADC_3bit_0/comp_p_6/vinn 0.19732f
C161 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin uo_out[2] 0.00138f
C162 uio_in[1] uio_in[0] 0.03102f
C163 flashADC_3bit_0/comp_p_1/out_left uio_out[0] 0
C164 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin -0
C165 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin 0
C166 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin uo_out[1] 0.00282f
C167 uo_out[7] uo_out[5] 0.00111f
C168 VDPWR uo_out[7] 1.68424f
C169 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A uo_out[0] 0
C170 uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B 0
C171 flashADC_3bit_0/comp_p_2/out_left VDPWR 0.14457f
C172 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VDPWR 0.02718f
C173 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in uo_out[1] 0.00492f
C174 uio_oe[5] VDPWR 0
C175 VDPWR uo_out[5] 1.25716f
C176 VDPWR uo_out[1] 0.017f
C177 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_4/latch_right -0.02778f
C178 uio_in[7] uio_in[6] 0.03102f
C179 uio_in[5] VDPWR 0
C180 ua[1] ua[0] 4.5498f
C181 flashADC_3bit_0/comp_p_6/vinn ua[0] 0
C182 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin uo_out[2] 0
C183 uo_out[7] uo_out[2] 0
C184 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in uo_out[2] 0
C185 VDPWR flashADC_3bit_0/comp_p_1/latch_right 0.22258f
C186 uo_out[5] uo_out[2] 0
C187 uo_out[2] uo_out[1] 2.07257f
C188 VDPWR uo_out[2] 0.08501f
C189 flashADC_3bit_0/comp_p_3/out_left VDPWR 0.18333f
C190 flashADC_3bit_0/comp_p_4/out_left flashADC_3bit_0/comp_p_5/vinn -0.00479f
C191 flashADC_3bit_0/comp_p_6/out_left VDPWR 0.26382f
C192 uio_oe[5] uio_oe[4] 0.03102f
C193 uo_out[3] uio_out[1] 0.00552f
C194 uo_out[6] uo_out[3] 0
C195 uio_oe[4] VDPWR 0
C196 uio_in[7] uo_out[0] 0.04843f
C197 uo_out[6] uo_out[4] 0
C198 flashADC_3bit_0/comp_p_6/vbias_p uio_out[1] 0.00692f
C199 uio_out[7] uio_oe[0] 0.03102f
C200 ui_in[3] ui_in[2] 0.03102f
C201 flashADC_3bit_0/vbias_generation_0/bias_n VDPWR 0.10568f
C202 flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_5/vinn -0.0296f
C203 uio_in[0] ui_in[7] 0.03102f
C204 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin uo_out[0] 0.00613f
C205 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.01661f
C206 uio_out[0] uo_out[7] 0.99679f
C207 ena clk 0.03102f
C208 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out VDPWR 1.28865f
C209 flashADC_3bit_0/comp_p_1/vinn uo_out[5] -0.0012f
C210 flashADC_3bit_0/comp_p_1/vinn VDPWR 1.17123f
C211 flashADC_3bit_0/comp_p_1/out_left uio_out[1] 0.03149f
C212 flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/comp_p_3/vinn -0.00404f
C213 flashADC_3bit_0/comp_p_3/vinn uo_out[5] -0.00952f
C214 uio_out[0] VDPWR 1.07221f
C215 uio_out[0] uo_out[5] 0
C216 VDPWR flashADC_3bit_0/comp_p_3/vinn 1.60219f
C217 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3] 0
C218 uio_out[3] uio_out[4] 0.03102f
C219 uio_in[6] uo_out[0] 0.01741f
C220 ua[7] ua[1] 0.01625f
C221 flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 VDPWR 0.03356f
C222 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G VDPWR 0.0124f
C223 uio_oe[3] VDPWR 0
C224 uio_in[4] uo_out[1] 0.01025f
C225 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 -0
C226 VDPWR flashADC_3bit_0/comp_p_0/vinn 1.85762f
C227 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in uo_out[0] 0.00561f
C228 uio_in[5] uio_in[4] 0.03102f
C229 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G uo_out[1] 0
C230 VDPWR flashADC_3bit_0/comp_p_6/latch_right 0.39269f
C231 uio_out[3] VDPWR 0
C232 ua[2] VGND 0.12712f
C233 ua[3] VGND 0.12712f
C234 ua[4] VGND 0.12712f
C235 ua[5] VGND 0.12712f
C236 ua[6] VGND 0.12712f
C237 ua[7] VGND 0.12842f
C238 ena VGND 0.07038f
C239 clk VGND 0.04288f
C240 rst_n VGND 0.04288f
C241 ui_in[0] VGND 0.04288f
C242 ui_in[1] VGND 0.04288f
C243 ui_in[2] VGND 0.04288f
C244 ui_in[3] VGND 0.04288f
C245 ui_in[4] VGND 0.04288f
C246 ui_in[5] VGND 0.04288f
C247 ui_in[6] VGND 0.04288f
C248 ui_in[7] VGND 0.04288f
C249 uio_in[0] VGND 0.04288f
C250 uio_in[1] VGND 0.04288f
C251 uio_in[2] VGND 0.04288f
C252 uio_in[3] VGND 0.03541f
C253 uio_in[4] VGND 0.03434f
C254 uio_in[5] VGND 0.0331f
C255 uio_in[6] VGND 0.0331f
C256 uio_in[7] VGND 0.0331f
C257 uio_out[2] VGND 0.04167f
C258 uio_out[3] VGND 0.04167f
C259 uio_out[4] VGND 0.04167f
C260 uio_out[5] VGND 0.04167f
C261 uio_out[6] VGND 0.04167f
C262 uio_out[7] VGND 0.04167f
C263 uio_oe[0] VGND 0.04176f
C264 uio_oe[1] VGND 0.04176f
C265 uio_oe[2] VGND 0.04167f
C266 uio_oe[3] VGND 0.04167f
C267 uio_oe[4] VGND 0.04167f
C268 uio_oe[5] VGND 0.04167f
C269 uio_oe[6] VGND 0.04167f
C270 uio_oe[7] VGND 0.06927f
C271 uo_out[2].n0 VGND 0.86264f
C272 uo_out[1].n0 VGND 0.90527f
C273 uio_out[1].t1 VGND 0.09868f
C274 uio_out[1].t0 VGND 0.09363f
C275 uio_out[1].n0 VGND 0.27936f
C276 uio_out[1].n1 VGND 2.99315f
C277 uio_out[1].n2 VGND 4.58739f
C278 flashADC_3bit_0/comp_p_6/out_left.t1 VGND 0.36236f
C279 flashADC_3bit_0/comp_p_6/out_left.n0 VGND 0.36336f
C280 flashADC_3bit_0/comp_p_6/out_left.t2 VGND 0.96524f
C281 flashADC_3bit_0/comp_p_6/out_left.n1 VGND 1.7499f
C282 flashADC_3bit_0/comp_p_6/out_left.t0 VGND 0.95737f
C283 flashADC_3bit_0/comp_p_6/out_left.n2 VGND 0.31727f
C284 flashADC_3bit_0/comp_p_6/out_left.n3 VGND 1.25549f
C285 uio_out[0].t0 VGND 0.12278f
C286 uio_out[0].t1 VGND 0.1294f
C287 uio_out[0].n0 VGND 0.36633f
C288 uio_out[0].n1 VGND 0.92016f
C289 uio_out[0].n2 VGND 5.10634f
C290 uo_out[7].t1 VGND 0.07979f
C291 uo_out[7].t0 VGND 0.07571f
C292 uo_out[7].n0 VGND 0.22588f
C293 uo_out[7].n1 VGND 4.90541f
C294 uo_out[7].n2 VGND 2.61036f
C295 flashADC_3bit_0/comp_p_4/out_left.t1 VGND 0.2858f
C296 flashADC_3bit_0/comp_p_4/out_left.n0 VGND 0.28659f
C297 flashADC_3bit_0/comp_p_4/out_left.t2 VGND 0.76131f
C298 flashADC_3bit_0/comp_p_4/out_left.n1 VGND 1.3802f
C299 flashADC_3bit_0/comp_p_4/out_left.t0 VGND 0.75511f
C300 flashADC_3bit_0/comp_p_4/out_left.n2 VGND 0.25024f
C301 flashADC_3bit_0/comp_p_4/out_left.n3 VGND 0.99025f
C302 uo_out[6].t0 VGND 0.10769f
C303 uo_out[6].t1 VGND 0.11349f
C304 uo_out[6].n0 VGND 0.3213f
C305 uo_out[6].n1 VGND 2.49197f
C306 uo_out[6].n2 VGND 0.38414f
C307 uo_out[6].n3 VGND 2.88453f
C308 flashADC_3bit_0/comp_p_3/out_left.t1 VGND 0.36236f
C309 flashADC_3bit_0/comp_p_3/out_left.n0 VGND 0.36336f
C310 flashADC_3bit_0/comp_p_3/out_left.t2 VGND 0.96524f
C311 flashADC_3bit_0/comp_p_3/out_left.n1 VGND 1.7499f
C312 flashADC_3bit_0/comp_p_3/out_left.t0 VGND 0.95737f
C313 flashADC_3bit_0/comp_p_3/out_left.n2 VGND 0.31727f
C314 flashADC_3bit_0/comp_p_3/out_left.n3 VGND 1.25549f
C315 flashADC_3bit_0/comp_p_3/latch_left.t0 VGND 1.27417f
C316 flashADC_3bit_0/comp_p_3/latch_left.t3 VGND 1.59739f
C317 flashADC_3bit_0/comp_p_3/latch_left.t2 VGND 1.48345f
C318 flashADC_3bit_0/comp_p_3/latch_left.n0 VGND 2.82036f
C319 flashADC_3bit_0/comp_p_3/latch_left.n1 VGND 1.81006f
C320 flashADC_3bit_0/comp_p_3/latch_left.t1 VGND 0.38095f
C321 flashADC_3bit_0/comp_p_3/latch_left.n2 VGND 1.62806f
C322 uo_out[5].t1 VGND 0.09276f
C323 uo_out[5].t0 VGND 0.08802f
C324 uo_out[5].n0 VGND 0.26072f
C325 uo_out[5].n1 VGND 0.05704f
C326 uo_out[5].n2 VGND 3.66875f
C327 uo_out[5].n3 VGND 2.20196f
C328 flashADC_3bit_0/comp_p_2/out_left.t1 VGND 0.27049f
C329 flashADC_3bit_0/comp_p_2/out_left.n0 VGND 0.27124f
C330 flashADC_3bit_0/comp_p_2/out_left.t2 VGND 0.72053f
C331 flashADC_3bit_0/comp_p_2/out_left.n1 VGND 1.30626f
C332 flashADC_3bit_0/comp_p_2/out_left.t0 VGND 0.71466f
C333 flashADC_3bit_0/comp_p_2/out_left.n2 VGND 0.23684f
C334 flashADC_3bit_0/comp_p_2/out_left.n3 VGND 0.9372f
C335 uo_out[4].t0 VGND 0.06216f
C336 uo_out[4].t1 VGND 0.06551f
C337 uo_out[4].n0 VGND 0.18546f
C338 uo_out[4].n1 VGND 2.98325f
C339 uo_out[4].n2 VGND 1.11497f
C340 flashADC_3bit_0/comp_p_0/latch_left.t0 VGND 1.01079f
C341 flashADC_3bit_0/comp_p_0/latch_left.t3 VGND 1.2672f
C342 flashADC_3bit_0/comp_p_0/latch_left.t2 VGND 1.17681f
C343 flashADC_3bit_0/comp_p_0/latch_left.n0 VGND 2.23738f
C344 flashADC_3bit_0/comp_p_0/latch_left.n1 VGND 1.43592f
C345 flashADC_3bit_0/comp_p_0/latch_left.t1 VGND 0.30221f
C346 flashADC_3bit_0/comp_p_0/latch_left.n2 VGND 1.29154f
C347 ua[0].t4 VGND 0.35499f
C348 ua[0].t5 VGND 0.35476f
C349 ua[0].n0 VGND 0.47665f
C350 ua[0].n1 VGND 0.37317f
C351 ua[0].t6 VGND 0.26383f
C352 ua[0].n2 VGND 0.4292f
C353 ua[0].t7 VGND 0.26349f
C354 ua[0].n3 VGND 0.42198f
C355 ua[0].n4 VGND 0.2f
C356 ua[0].t8 VGND 0.35499f
C357 ua[0].t9 VGND 0.35476f
C358 ua[0].n5 VGND 0.47665f
C359 ua[0].n6 VGND 0.37317f
C360 ua[0].t10 VGND 0.26383f
C361 ua[0].n7 VGND 0.4292f
C362 ua[0].t11 VGND 0.26349f
C363 ua[0].n8 VGND 0.42198f
C364 ua[0].n9 VGND 0.2f
C365 ua[0].n10 VGND 2.93699f
C366 ua[0].t16 VGND 0.35499f
C367 ua[0].t17 VGND 0.35476f
C368 ua[0].n11 VGND 0.47665f
C369 ua[0].n12 VGND 0.37317f
C370 ua[0].t18 VGND 0.26383f
C371 ua[0].n13 VGND 0.4292f
C372 ua[0].t19 VGND 0.26349f
C373 ua[0].n14 VGND 0.42198f
C374 ua[0].n15 VGND 0.2f
C375 ua[0].n16 VGND 1.89166f
C376 ua[0].n17 VGND 1.59712f
C377 ua[0].t24 VGND 0.35499f
C378 ua[0].t25 VGND 0.35476f
C379 ua[0].n18 VGND 0.47665f
C380 ua[0].n19 VGND 0.37317f
C381 ua[0].t26 VGND 0.26383f
C382 ua[0].n20 VGND 0.4292f
C383 ua[0].t27 VGND 0.26349f
C384 ua[0].n21 VGND 0.42198f
C385 ua[0].n22 VGND 0.2f
C386 ua[0].t0 VGND 0.35499f
C387 ua[0].t1 VGND 0.35476f
C388 ua[0].n23 VGND 0.47665f
C389 ua[0].n24 VGND 0.37317f
C390 ua[0].t2 VGND 0.26383f
C391 ua[0].n25 VGND 0.4292f
C392 ua[0].t3 VGND 0.26349f
C393 ua[0].n26 VGND 0.42198f
C394 ua[0].n27 VGND 0.19355f
C395 ua[0].n28 VGND 0.90835f
C396 ua[0].t12 VGND 0.35499f
C397 ua[0].t13 VGND 0.35476f
C398 ua[0].n29 VGND 0.47665f
C399 ua[0].n30 VGND 0.37317f
C400 ua[0].t14 VGND 0.26383f
C401 ua[0].n31 VGND 0.4292f
C402 ua[0].t15 VGND 0.26349f
C403 ua[0].n32 VGND 0.42198f
C404 ua[0].n33 VGND 0.19893f
C405 ua[0].n34 VGND 0.20405f
C406 ua[0].n35 VGND 3.03157f
C407 ua[0].t20 VGND 0.35499f
C408 ua[0].t21 VGND 0.35476f
C409 ua[0].n36 VGND 0.47665f
C410 ua[0].n37 VGND 0.37317f
C411 ua[0].t22 VGND 0.26383f
C412 ua[0].n38 VGND 0.4292f
C413 ua[0].t23 VGND 0.26349f
C414 ua[0].n39 VGND 0.42198f
C415 ua[0].n40 VGND 0.19539f
C416 ua[0].n41 VGND 0.2648f
C417 ua[0].n42 VGND 2.35755f
C418 ua[0].n43 VGND 2.16931f
C419 ua[0].n44 VGND 1.15796f
C420 ua[0].n45 VGND 0.80821f
C421 uo_out[3].t1 VGND 0.06421f
C422 uo_out[3].t0 VGND 0.06093f
C423 uo_out[3].n0 VGND 0.18004f
C424 uo_out[3].n1 VGND 0.04119f
C425 uo_out[3].n2 VGND 1.07213f
C426 uo_out[3].n3 VGND 1.08672f
C427 flashADC_3bit_0/comp_p_1/out_left.t1 VGND 0.36236f
C428 flashADC_3bit_0/comp_p_1/out_left.n0 VGND 0.36336f
C429 flashADC_3bit_0/comp_p_1/out_left.t2 VGND 0.96524f
C430 flashADC_3bit_0/comp_p_1/out_left.n1 VGND 1.7499f
C431 flashADC_3bit_0/comp_p_1/out_left.t0 VGND 0.95737f
C432 flashADC_3bit_0/comp_p_1/out_left.n2 VGND 0.31727f
C433 flashADC_3bit_0/comp_p_1/out_left.n3 VGND 1.25549f
C434 ua[1].n0 VGND 0.50626f
C435 ua[1].n1 VGND 2.58175f
C436 VDPWR.n0 VGND 0.44704f
C437 VDPWR.n1 VGND 0.65278f
C438 VDPWR.n2 VGND 1.31241f
C439 VDPWR.n3 VGND 13.2291f
C440 VDPWR.n4 VGND 0.00781f
C441 VDPWR.n5 VGND 0.01558f
C442 VDPWR.n6 VGND 0.12532f
C443 VDPWR.n7 VGND 0.0152f
C444 VDPWR.n8 VGND 0.11439f
C445 VDPWR.n9 VGND 0.01558f
C446 VDPWR.n10 VGND 0.01558f
C447 VDPWR.n11 VGND 0.00544f
C448 VDPWR.n12 VGND 0.00781f
C449 VDPWR.n13 VGND 0.11439f
C450 VDPWR.n14 VGND 0.01011f
C451 VDPWR.n15 VGND 0.01011f
C452 VDPWR.n16 VGND 0.01011f
C453 VDPWR.n17 VGND 0.01025f
C454 VDPWR.n18 VGND 0.00977f
C455 VDPWR.n19 VGND 0.00977f
C456 VDPWR.n20 VGND 0.00977f
C457 VDPWR.n21 VGND 0.11439f
C458 VDPWR.n22 VGND 0.11439f
C459 VDPWR.n23 VGND 0.00977f
C460 VDPWR.n24 VGND 0.01025f
C461 VDPWR.n25 VGND 0.00977f
C462 VDPWR.n26 VGND 0.0152f
C463 VDPWR.n27 VGND 0.0152f
C464 VDPWR.n28 VGND 0.11439f
C465 VDPWR.n29 VGND 0.01558f
C466 VDPWR.n30 VGND 0.01558f
C467 VDPWR.n31 VGND 0.00544f
C468 VDPWR.n32 VGND 0.00781f
C469 VDPWR.n33 VGND 0.12532f
C470 VDPWR.n34 VGND 0.01558f
C471 VDPWR.n35 VGND 0.01558f
C472 VDPWR.n36 VGND 0.07278f
C473 VDPWR.n37 VGND 0.04324f
C474 VDPWR.n38 VGND 0.14024f
C475 VDPWR.n39 VGND 0.00766f
C476 VDPWR.n40 VGND 0.00781f
C477 VDPWR.n42 VGND 0.09985f
C478 VDPWR.n43 VGND 0.0152f
C479 VDPWR.n44 VGND 0.01519f
C480 VDPWR.n45 VGND 0.0152f
C481 VDPWR.n46 VGND 0.09485f
C482 VDPWR.n47 VGND 0.09485f
C483 VDPWR.n48 VGND 0.0152f
C484 VDPWR.n49 VGND 0.0152f
C485 VDPWR.n50 VGND 0.01519f
C486 VDPWR.n51 VGND 0.0152f
C487 VDPWR.n52 VGND 0.47712f
C488 VDPWR.n53 VGND 0.47712f
C489 VDPWR.n54 VGND 0.01011f
C490 VDPWR.n55 VGND 0.11439f
C491 VDPWR.n56 VGND 0.01011f
C492 VDPWR.n57 VGND 0.01011f
C493 VDPWR.n58 VGND 0.01025f
C494 VDPWR.n59 VGND 0.01025f
C495 VDPWR.n60 VGND 0.00977f
C496 VDPWR.n61 VGND 0.00975f
C497 VDPWR.n62 VGND 0.07278f
C498 VDPWR.n63 VGND 0.04349f
C499 VDPWR.n64 VGND 0.11496f
C500 VDPWR.n65 VGND 0.12132f
C501 VDPWR.n66 VGND 0.00232f
C502 VDPWR.n67 VGND 0.00234f
C503 VDPWR.n68 VGND 0.00464f
C504 VDPWR.n69 VGND 0.11439f
C505 VDPWR.n70 VGND 0.00464f
C506 VDPWR.n71 VGND 0.00977f
C507 VDPWR.n72 VGND 0.0152f
C508 VDPWR.n73 VGND 0.0152f
C509 VDPWR.n74 VGND 0.09557f
C510 VDPWR.n75 VGND 0.09557f
C511 VDPWR.n76 VGND 0.0152f
C512 VDPWR.n77 VGND 0.0152f
C513 VDPWR.n78 VGND 0.01519f
C514 VDPWR.n79 VGND 0.0152f
C515 VDPWR.n80 VGND 0.09485f
C516 VDPWR.n81 VGND 0.09485f
C517 VDPWR.n82 VGND 0.0152f
C518 VDPWR.n83 VGND 0.01558f
C519 VDPWR.n85 VGND 0.09985f
C520 VDPWR.n86 VGND 0.01519f
C521 VDPWR.n87 VGND 0.00544f
C522 VDPWR.n88 VGND 0.04324f
C523 VDPWR.n89 VGND 0.07278f
C524 VDPWR.n90 VGND 1.12518f
C525 VDPWR.n91 VGND 1.73918f
C526 VDPWR.n92 VGND 0.51635f
C527 VDPWR.n93 VGND 0.36214f
C528 VDPWR.n94 VGND 0.01419f
C529 VDPWR.n95 VGND 0.08043f
C530 VDPWR.n96 VGND 0.36214f
C531 VDPWR.n97 VGND 0.39067f
C532 VDPWR.n98 VGND 0.01752f
C533 VDPWR.n99 VGND 0.21055f
C534 VDPWR.n100 VGND 0.0317f
C535 VDPWR.n101 VGND 0.03582f
C536 VDPWR.n102 VGND 2.23986f
C537 VDPWR.n103 VGND 0.03179f
C538 VDPWR.n104 VGND 0.03179f
C539 VDPWR.n105 VGND 0.40354f
C540 VDPWR.n106 VGND 0.0317f
C541 VDPWR.n107 VGND 0.03582f
C542 VDPWR.n108 VGND 0.11569f
C543 VDPWR.n109 VGND -0.08122f
C544 VDPWR.n110 VGND 0.01752f
C545 VDPWR.n111 VGND 0.03582f
C546 VDPWR.n112 VGND 0.02935f
C547 VDPWR.n113 VGND 0.50329f
C548 VDPWR.n114 VGND 0.03179f
C549 VDPWR.n115 VGND 2.18998f
C550 VDPWR.n116 VGND 0.03179f
C551 VDPWR.n117 VGND 0.10703f
C552 VDPWR.n118 VGND 0.20877f
C553 VDPWR.n119 VGND 0.65864f
C554 VDPWR.n120 VGND 0.04105f
C555 VDPWR.n121 VGND 0.04105f
C556 VDPWR.n122 VGND 2.45523f
C557 VDPWR.n123 VGND 0.04105f
C558 VDPWR.n124 VGND 0.04105f
C559 VDPWR.n125 VGND 0.02935f
C560 VDPWR.n126 VGND 0.03582f
C561 VDPWR.n127 VGND 0.20877f
C562 VDPWR.n128 VGND 0.65864f
C563 VDPWR.n129 VGND 0.10703f
C564 VDPWR.n130 VGND 0.10628f
C565 VDPWR.n131 VGND 0.11466f
C566 VDPWR.n132 VGND 0.37096f
C567 VDPWR.n133 VGND 0.04082f
C568 VDPWR.n134 VGND 0.04097f
C569 VDPWR.n135 VGND 0.67433f
C570 VDPWR.n136 VGND 0.22059f
C571 VDPWR.n137 VGND 2.55724f
C572 VDPWR.n138 VGND 0.04097f
C573 VDPWR.n139 VGND 0.04097f
C574 VDPWR.n140 VGND 0.10628f
C575 VDPWR.n141 VGND 0.11466f
C576 VDPWR.n142 VGND 0.01489f
C577 VDPWR.n143 VGND 0.21937f
C578 VDPWR.n144 VGND 2.55724f
C579 VDPWR.n145 VGND 0.04904f
C580 VDPWR.n146 VGND 0.04097f
C581 VDPWR.n147 VGND 0.04097f
C582 VDPWR.n148 VGND 0.67433f
C583 VDPWR.n149 VGND 0.01489f
C584 VDPWR.n150 VGND 0.21937f
C585 VDPWR.n151 VGND 0.04884f
C586 VDPWR.n152 VGND 0.04082f
C587 VDPWR.n153 VGND 1.79778f
C588 VDPWR.n154 VGND 0.04096f
C589 VDPWR.n155 VGND 0.04096f
C590 VDPWR.n156 VGND 2.53231f
C591 VDPWR.n157 VGND 0.04884f
C592 VDPWR.n158 VGND 0.04082f
C593 VDPWR.n159 VGND 0.21937f
C594 VDPWR.n160 VGND 0.01489f
C595 VDPWR.n161 VGND 0.22059f
C596 VDPWR.n162 VGND 2.56858f
C597 VDPWR.n163 VGND 0.04097f
C598 VDPWR.n164 VGND 0.04173f
C599 VDPWR.n165 VGND 0.04105f
C600 VDPWR.n166 VGND 0.04105f
C601 VDPWR.n167 VGND 0.1065f
C602 VDPWR.n168 VGND 0.04173f
C603 VDPWR.n169 VGND 0.35958f
C604 VDPWR.n170 VGND -0.08122f
C605 VDPWR.n171 VGND 0.03582f
C606 VDPWR.n172 VGND 0.00664f
C607 VDPWR.n173 VGND 0.03179f
C608 VDPWR.n174 VGND 0.10405f
C609 VDPWR.n175 VGND 0.00664f
C610 VDPWR.n176 VGND 0.65864f
C611 VDPWR.n177 VGND 0.20877f
C612 VDPWR.n178 VGND 0.0317f
C613 VDPWR.n179 VGND 0.03179f
C614 VDPWR.n180 VGND 0.02935f
C615 VDPWR.n181 VGND 0.01752f
C616 VDPWR.n182 VGND 0.6806f
C617 VDPWR.n183 VGND 0.39067f
C618 VDPWR.n184 VGND 0.01752f
C619 VDPWR.n185 VGND 0.21055f
C620 VDPWR.n186 VGND 0.0317f
C621 VDPWR.n187 VGND 0.0317f
C622 VDPWR.n188 VGND 0.10405f
C623 VDPWR.n189 VGND 0.67433f
C624 VDPWR.n190 VGND 0.37096f
C625 VDPWR.n191 VGND 0.0058f
C626 VDPWR.n192 VGND 0.10703f
C627 VDPWR.n193 VGND 0.04173f
C628 VDPWR.n194 VGND 0.01923f
C629 VDPWR.n195 VGND 0.03179f
C630 VDPWR.n196 VGND 0.35958f
C631 VDPWR.n197 VGND 0.65864f
C632 VDPWR.n198 VGND 0.02935f
C633 VDPWR.n199 VGND 0.20877f
C634 VDPWR.n200 VGND 2.08343f
C635 VDPWR.n201 VGND 2.45523f
C636 VDPWR.n202 VGND 0.03582f
C637 VDPWR.n203 VGND 0.03179f
C638 VDPWR.n204 VGND 0.11157f
C639 VDPWR.n205 VGND -0.08122f
C640 VDPWR.n206 VGND 0.04105f
C641 VDPWR.n207 VGND 0.04082f
C642 VDPWR.n208 VGND 0.01489f
C643 VDPWR.n209 VGND 0.00664f
C644 VDPWR.n210 VGND 0.00664f
C645 VDPWR.n211 VGND 0.04082f
C646 VDPWR.n212 VGND 0.01489f
C647 VDPWR.n213 VGND 2.23986f
C648 VDPWR.n214 VGND 2.18998f
C649 VDPWR.n215 VGND 0.04105f
C650 VDPWR.n216 VGND 0.10628f
C651 VDPWR.n217 VGND 0.11466f
C652 VDPWR.n218 VGND 0.11569f
C653 VDPWR.n219 VGND 0.1065f
C654 VDPWR.n220 VGND 0.03179f
C655 VDPWR.n221 VGND 0.03582f
C656 VDPWR.n222 VGND 0.03179f
C657 VDPWR.n223 VGND 0.02931f
C658 VDPWR.n224 VGND 0.01419f
C659 VDPWR.n225 VGND 0.02338f
C660 VDPWR.n226 VGND 0.01419f
C661 VDPWR.n227 VGND 0.02931f
C662 VDPWR.n228 VGND 0.21055f
C663 VDPWR.n229 VGND 0.03582f
C664 VDPWR.n230 VGND 0.03179f
C665 VDPWR.n231 VGND 0.0317f
C666 VDPWR.n232 VGND 0.03179f
C667 VDPWR.n233 VGND 0.11157f
C668 VDPWR.n234 VGND 0.01923f
C669 VDPWR.n235 VGND 0.10703f
C670 VDPWR.n236 VGND 0.10628f
C671 VDPWR.n237 VGND 0.11466f
C672 VDPWR.n238 VGND 0.11569f
C673 VDPWR.n239 VGND 0.0058f
C674 VDPWR.n240 VGND 0.37096f
C675 VDPWR.n241 VGND 0.04173f
C676 VDPWR.n242 VGND 1.81138f
C677 VDPWR.n243 VGND 0.40354f
C678 VDPWR.n244 VGND 0.04097f
C679 VDPWR.n245 VGND 0.03765f
C680 VDPWR.n246 VGND 0.04082f
C681 VDPWR.n247 VGND 0.03765f
C682 VDPWR.n248 VGND 0.04096f
C683 VDPWR.n249 VGND 0.50329f
C684 VDPWR.n250 VGND 0.04096f
C685 VDPWR.n251 VGND 0.03765f
C686 VDPWR.n252 VGND 0.04082f
C687 VDPWR.n253 VGND 0.03765f
C688 VDPWR.n254 VGND 0.22059f
C689 VDPWR.n255 VGND 0.04904f
C690 VDPWR.n256 VGND 2.6774f
C691 VDPWR.n257 VGND 0.04096f
C692 VDPWR.n258 VGND 0.04096f
C693 VDPWR.n259 VGND 0.03765f
C694 VDPWR.n260 VGND 0.04082f
C695 VDPWR.n261 VGND 0.01489f
C696 VDPWR.n262 VGND 0.01489f
C697 VDPWR.n263 VGND 0.04082f
C698 VDPWR.n264 VGND 0.03765f
C699 VDPWR.n265 VGND 0.21937f
C700 VDPWR.n266 VGND 0.04884f
C701 VDPWR.n267 VGND 2.67513f
C702 VDPWR.n268 VGND 0.04884f
C703 VDPWR.n269 VGND 0.04096f
C704 VDPWR.n270 VGND 0.04082f
C705 VDPWR.n271 VGND 0.01489f
C706 VDPWR.n272 VGND 0.04082f
C707 VDPWR.n273 VGND 0.04096f
C708 VDPWR.n274 VGND 0.03765f
C709 VDPWR.n275 VGND 0.04082f
C710 VDPWR.n276 VGND 0.03765f
C711 VDPWR.n277 VGND 0.02931f
C712 VDPWR.n278 VGND 0.21055f
C713 VDPWR.n279 VGND 0.0058f
C714 VDPWR.n280 VGND 0.04173f
C715 VDPWR.n281 VGND 1.81138f
C716 VDPWR.n282 VGND 0.04173f
C717 VDPWR.n283 VGND 0.37096f
C718 VDPWR.n284 VGND 0.67433f
C719 VDPWR.n285 VGND 0.22059f
C720 VDPWR.n286 VGND 0.04904f
C721 VDPWR.n287 VGND 2.08116f
C722 VDPWR.n288 VGND 0.04904f
C723 VDPWR.n289 VGND 0.04097f
C724 VDPWR.n290 VGND 0.0058f
C725 VDPWR.n291 VGND 0.11569f
C726 VDPWR.n292 VGND 0.1065f
C727 VDPWR.n293 VGND 0.0317f
C728 VDPWR.n294 VGND 0.00664f
C729 VDPWR.n295 VGND 0.00664f
C730 VDPWR.n296 VGND 0.10405f
C731 VDPWR.n297 VGND -0.08122f
C732 VDPWR.n298 VGND 0.11157f
C733 VDPWR.n299 VGND 0.01923f
C734 VDPWR.n300 VGND 0.35958f
C735 VDPWR.n301 VGND 0.04173f
C736 VDPWR.n302 VGND 1.79778f
C737 VDPWR.n303 VGND 0.04173f
C738 VDPWR.n304 VGND 0.35958f
C739 VDPWR.n305 VGND 0.01923f
C740 VDPWR.n306 VGND 0.11157f
C741 VDPWR.n307 VGND 0.03179f
C742 VDPWR.n308 VGND 2.53231f
C743 VDPWR.n309 VGND 0.03179f
C744 VDPWR.n310 VGND 0.0317f
C745 VDPWR.n311 VGND 0.00664f
C746 VDPWR.n312 VGND 0.00664f
C747 VDPWR.n313 VGND 0.10405f
C748 VDPWR.n314 VGND 0.1065f
C749 VDPWR.n315 VGND 0.03179f
C750 VDPWR.n316 VGND 2.56858f
C751 VDPWR.n317 VGND 0.03179f
C752 VDPWR.n318 VGND 0.02931f
C753 VDPWR.n319 VGND 0.01419f
C754 VDPWR.n320 VGND 0.02338f
C755 VDPWR.n321 VGND 0.6806f
C756 VDPWR.n322 VGND 0.51622f
C757 VDPWR.n323 VGND 3.01936f
C758 VDPWR.n324 VGND 0.1851f
C759 VDPWR.n325 VGND 0.14048f
C760 VDPWR.n326 VGND 0.1216f
C761 VDPWR.n327 VGND 0.2109f
C762 VDPWR.n328 VGND 0.40426f
C763 VDPWR.n329 VGND 0.56037f
C764 VDPWR.n330 VGND 0.01752f
C765 VDPWR.n331 VGND 0.21055f
C766 VDPWR.n332 VGND 0.0317f
C767 VDPWR.n333 VGND 0.03582f
C768 VDPWR.n334 VGND 1.11993f
C769 VDPWR.n335 VGND 0.03179f
C770 VDPWR.n336 VGND 0.04097f
C771 VDPWR.n337 VGND 0.90569f
C772 VDPWR.n338 VGND 0.04082f
C773 VDPWR.n339 VGND 1.38646f
C774 VDPWR.n340 VGND 0.98179f
C775 VDPWR.n341 VGND 0.11569f
C776 VDPWR.n342 VGND 0.67433f
C777 VDPWR.n343 VGND 0.04105f
C778 VDPWR.n344 VGND 0.04173f
C779 VDPWR.n345 VGND 0.10628f
C780 VDPWR.n346 VGND 0.25164f
C781 VDPWR.n347 VGND 0.03179f
C782 VDPWR.n348 VGND 0.03582f
C783 VDPWR.n349 VGND 0.21937f
C784 VDPWR.n350 VGND 0.04082f
C785 VDPWR.n351 VGND 0.22059f
C786 VDPWR.n352 VGND 0.03765f
C787 VDPWR.n353 VGND 0.11466f
C788 VDPWR.n354 VGND 0.01489f
C789 VDPWR.n355 VGND 0.01489f
C790 VDPWR.n356 VGND 0.04082f
C791 VDPWR.n357 VGND 0.03765f
C792 VDPWR.n358 VGND 0.04096f
C793 VDPWR.n359 VGND 1.27862f
C794 VDPWR.n360 VGND 0.04097f
C795 VDPWR.n361 VGND 0.04097f
C796 VDPWR.n362 VGND 0.67433f
C797 VDPWR.n363 VGND 0.01489f
C798 VDPWR.n364 VGND 0.21937f
C799 VDPWR.n365 VGND 0.98231f
C800 VDPWR.n366 VGND 0.04082f
C801 VDPWR.n367 VGND 0.89889f
C802 VDPWR.n368 VGND 0.04096f
C803 VDPWR.n369 VGND 0.03179f
C804 VDPWR.n370 VGND 1.09499f
C805 VDPWR.n371 VGND 1.33585f
C806 VDPWR.n372 VGND 0.03582f
C807 VDPWR.n373 VGND 0.0317f
C808 VDPWR.n374 VGND 0.20877f
C809 VDPWR.n375 VGND 0.00664f
C810 VDPWR.n376 VGND 0.21055f
C811 VDPWR.n377 VGND 0.03582f
C812 VDPWR.n378 VGND 0.04082f
C813 VDPWR.n379 VGND 0.01489f
C814 VDPWR.n380 VGND 1.11993f
C815 VDPWR.n381 VGND 0.00664f
C816 VDPWR.n382 VGND 0.0317f
C817 VDPWR.n383 VGND 0.03179f
C818 VDPWR.n384 VGND 0.04105f
C819 VDPWR.n385 VGND 0.04105f
C820 VDPWR.n386 VGND 0.1065f
C821 VDPWR.n387 VGND 0.65864f
C822 VDPWR.n388 VGND 0.04173f
C823 VDPWR.n389 VGND 0.35958f
C824 VDPWR.n390 VGND 0.10405f
C825 VDPWR.n391 VGND -0.08122f
C826 VDPWR.n392 VGND 0.11157f
C827 VDPWR.n393 VGND 0.01923f
C828 VDPWR.n394 VGND 0.10703f
C829 VDPWR.n395 VGND 0.10628f
C830 VDPWR.n396 VGND 0.11466f
C831 VDPWR.n397 VGND 0.11569f
C832 VDPWR.n398 VGND 0.0058f
C833 VDPWR.n399 VGND 0.37096f
C834 VDPWR.n400 VGND 0.04173f
C835 VDPWR.n401 VGND 0.90569f
C836 VDPWR.n402 VGND 0.20177f
C837 VDPWR.n403 VGND 1.28429f
C838 VDPWR.n404 VGND 0.03179f
C839 VDPWR.n405 VGND 0.02931f
C840 VDPWR.n406 VGND 0.73719f
C841 VDPWR.n407 VGND 0.79353f
C842 VDPWR.n408 VGND 1.76274f
C843 VDPWR.n409 VGND 0.28982f
C844 VDPWR.n410 VGND 0.40401f
C845 VDPWR.n411 VGND 0.56037f
C846 VDPWR.n412 VGND 0.04337f
C847 VDPWR.n413 VGND 0.01419f
C848 VDPWR.n414 VGND 0.01752f
C849 VDPWR.n415 VGND 0.02935f
C850 VDPWR.n416 VGND 0.03179f
C851 VDPWR.n417 VGND 1.26615f
C852 VDPWR.n418 VGND 0.25164f
C853 VDPWR.n419 VGND 0.04096f
C854 VDPWR.n420 VGND 0.03765f
C855 VDPWR.n421 VGND 0.04082f
C856 VDPWR.n422 VGND 0.03765f
C857 VDPWR.n423 VGND 0.22059f
C858 VDPWR.n424 VGND 0.04904f
C859 VDPWR.n425 VGND 1.3387f
C860 VDPWR.n426 VGND 0.89889f
C861 VDPWR.n427 VGND 1.22761f
C862 VDPWR.n428 VGND 1.33757f
C863 VDPWR.n429 VGND 0.04884f
C864 VDPWR.n430 VGND 0.04096f
C865 VDPWR.n431 VGND 0.10703f
C866 VDPWR.n432 VGND 0.1065f
C867 VDPWR.n433 VGND 0.0317f
C868 VDPWR.n434 VGND 0.00664f
C869 VDPWR.n435 VGND 0.00664f
C870 VDPWR.n436 VGND 0.10405f
C871 VDPWR.n437 VGND -0.08122f
C872 VDPWR.n438 VGND 0.11157f
C873 VDPWR.n439 VGND 0.01923f
C874 VDPWR.n440 VGND 0.35958f
C875 VDPWR.n441 VGND 0.65864f
C876 VDPWR.n442 VGND 0.20877f
C877 VDPWR.n443 VGND 0.02935f
C878 VDPWR.n444 VGND 0.03179f
C879 VDPWR.n445 VGND 1.26615f
C880 VDPWR.n446 VGND 1.09499f
C881 VDPWR.n447 VGND 0.04105f
C882 VDPWR.n448 VGND 0.04173f
C883 VDPWR.n449 VGND 0.37096f
C884 VDPWR.n450 VGND 0.0058f
C885 VDPWR.n451 VGND 0.04097f
C886 VDPWR.n452 VGND 0.20177f
C887 VDPWR.n453 VGND 1.28429f
C888 VDPWR.n454 VGND 0.03179f
C889 VDPWR.n455 VGND 0.02931f
C890 VDPWR.n456 VGND 0.01419f
C891 VDPWR.n457 VGND 0.04337f
C892 VDPWR.n458 VGND 0.73719f
C893 VDPWR.n459 VGND 0.79353f
C894 VDPWR.n460 VGND 2.00287f
C895 VDPWR.n461 VGND 0.15605f
C896 VDPWR.n462 VGND 1.14311f
C897 VDPWR.n463 VGND 1.99909f
C898 VDPWR.n464 VGND 1.16102f
C899 VDPWR.n465 VGND 2.69599f
C900 VDPWR.n466 VGND 3.54107f
C901 VDPWR.n467 VGND 3.63065f
C902 VDPWR.n468 VGND 3.91276f
C903 VDPWR.n469 VGND 0.00544f
C904 VDPWR.n470 VGND 0.10818f
C905 VDPWR.n471 VGND 0.00781f
C906 VDPWR.n472 VGND 0.01558f
C907 VDPWR.n473 VGND 0.01558f
C908 VDPWR.n474 VGND 0.77318f
C909 VDPWR.n475 VGND 0.0152f
C910 VDPWR.n476 VGND 0.77318f
C911 VDPWR.n477 VGND 0.0152f
C912 VDPWR.n478 VGND 0.0152f
C913 VDPWR.n479 VGND 0.01558f
C914 VDPWR.n480 VGND 0.01558f
C915 VDPWR.n481 VGND 0.01519f
C916 VDPWR.n482 VGND 0.00781f
C917 VDPWR.n483 VGND 0.01558f
C918 VDPWR.n484 VGND 0.01558f
C919 VDPWR.n485 VGND 0.77318f
C920 VDPWR.n486 VGND 0.0152f
C921 VDPWR.n487 VGND 0.0152f
C922 VDPWR.n488 VGND 0.0152f
C923 VDPWR.n489 VGND 0.77318f
C924 VDPWR.n490 VGND 0.01558f
C925 VDPWR.n491 VGND 0.01558f
C926 VDPWR.n492 VGND 0.00781f
C927 VDPWR.n493 VGND 0.0152f
C928 VDPWR.n494 VGND 0.01519f
C929 VDPWR.n495 VGND 0.0152f
C930 VDPWR.n496 VGND 1.19908f
C931 VDPWR.n497 VGND 0.0152f
C932 VDPWR.n498 VGND 0.01519f
C933 VDPWR.n499 VGND 0.00544f
C934 VDPWR.n500 VGND 0.10818f
C935 VDPWR.n501 VGND 0.02419f
C936 VDPWR.n502 VGND 0.00544f
C937 VDPWR.n503 VGND 0.00781f
C938 VDPWR.n504 VGND 0.0152f
C939 VDPWR.n505 VGND 0.0152f
C940 VDPWR.n506 VGND 1.19908f
C941 VDPWR.n507 VGND 0.0152f
C942 VDPWR.n508 VGND 0.01519f
C943 VDPWR.n509 VGND 0.00544f
C944 VDPWR.n510 VGND 0.12229f
C945 VDPWR.n511 VGND 0.66459f
C946 VDPWR.n512 VGND 1.18891f
C947 VDPWR.n513 VGND 0.65638f
C948 VDPWR.n514 VGND 3.6595f
C949 VDPWR.n515 VGND 1.75044f
C950 VDPWR.n516 VGND 0.78025f
C951 VDPWR.n517 VGND 0.00544f
C952 VDPWR.n518 VGND 0.10818f
C953 VDPWR.n519 VGND 0.00781f
C954 VDPWR.n520 VGND 0.01558f
C955 VDPWR.n521 VGND 0.01558f
C956 VDPWR.n522 VGND 0.77318f
C957 VDPWR.n523 VGND 0.0152f
C958 VDPWR.n524 VGND 0.77318f
C959 VDPWR.n525 VGND 0.0152f
C960 VDPWR.n526 VGND 0.0152f
C961 VDPWR.n527 VGND 0.01558f
C962 VDPWR.n528 VGND 0.01558f
C963 VDPWR.n529 VGND 0.01519f
C964 VDPWR.n530 VGND 0.00781f
C965 VDPWR.n531 VGND 0.01558f
C966 VDPWR.n532 VGND 0.01558f
C967 VDPWR.n533 VGND 0.77318f
C968 VDPWR.n534 VGND 0.0152f
C969 VDPWR.n535 VGND 0.0152f
C970 VDPWR.n536 VGND 0.0152f
C971 VDPWR.n537 VGND 0.77318f
C972 VDPWR.n538 VGND 0.01558f
C973 VDPWR.n539 VGND 0.01558f
C974 VDPWR.n540 VGND 0.00781f
C975 VDPWR.n541 VGND 0.0152f
C976 VDPWR.n542 VGND 0.01519f
C977 VDPWR.n543 VGND 0.0152f
C978 VDPWR.n544 VGND 1.19908f
C979 VDPWR.n545 VGND 0.0152f
C980 VDPWR.n546 VGND 0.01519f
C981 VDPWR.n547 VGND 0.00544f
C982 VDPWR.n548 VGND 0.10818f
C983 VDPWR.n549 VGND 0.02419f
C984 VDPWR.n550 VGND 0.00544f
C985 VDPWR.n551 VGND 0.00781f
C986 VDPWR.n552 VGND 0.0152f
C987 VDPWR.n553 VGND 0.0152f
C988 VDPWR.n554 VGND 1.19908f
C989 VDPWR.n555 VGND 0.0152f
C990 VDPWR.n556 VGND 0.01519f
C991 VDPWR.n557 VGND 0.00544f
C992 VDPWR.n558 VGND 0.12229f
C993 VDPWR.n559 VGND 0.66576f
C994 VDPWR.n560 VGND 0.71657f
C995 VDPWR.n561 VGND 1.8337f
C996 VDPWR.n562 VGND 3.11532f
C997 VDPWR.n563 VGND 0.59065f
C998 VDPWR.n564 VGND 0.08969f
C999 VDPWR.n565 VGND 0.21386f
C1000 VDPWR.n566 VGND 1.42105f
C1001 VDPWR.n567 VGND 0.55544f
C1002 VDPWR.n568 VGND 0.4649f
C1003 VDPWR.n569 VGND 0.46453f
C1004 VDPWR.n570 VGND 0.58691f
C1005 VDPWR.n571 VGND 0.01752f
C1006 VDPWR.n572 VGND 0.21055f
C1007 VDPWR.n573 VGND 0.0317f
C1008 VDPWR.n574 VGND 0.03582f
C1009 VDPWR.n575 VGND 1.11993f
C1010 VDPWR.n576 VGND 0.03179f
C1011 VDPWR.n577 VGND 0.04097f
C1012 VDPWR.n578 VGND 0.90569f
C1013 VDPWR.n579 VGND 0.04082f
C1014 VDPWR.n580 VGND 1.38646f
C1015 VDPWR.n581 VGND 0.98179f
C1016 VDPWR.n582 VGND 0.11569f
C1017 VDPWR.n583 VGND 0.67433f
C1018 VDPWR.n584 VGND 0.04105f
C1019 VDPWR.n585 VGND 0.04173f
C1020 VDPWR.n586 VGND -0.08122f
C1021 VDPWR.n587 VGND 0.25164f
C1022 VDPWR.n588 VGND 0.1065f
C1023 VDPWR.n589 VGND 0.10405f
C1024 VDPWR.n590 VGND 0.00664f
C1025 VDPWR.n591 VGND 0.00664f
C1026 VDPWR.n592 VGND 0.0317f
C1027 VDPWR.n593 VGND 0.03179f
C1028 VDPWR.n594 VGND 0.03582f
C1029 VDPWR.n595 VGND 0.21937f
C1030 VDPWR.n596 VGND 0.10628f
C1031 VDPWR.n597 VGND 0.04082f
C1032 VDPWR.n598 VGND 0.11466f
C1033 VDPWR.n599 VGND 0.01489f
C1034 VDPWR.n600 VGND 0.01489f
C1035 VDPWR.n601 VGND 0.22059f
C1036 VDPWR.n602 VGND 0.03765f
C1037 VDPWR.n603 VGND 0.04082f
C1038 VDPWR.n604 VGND 0.03765f
C1039 VDPWR.n605 VGND 0.04096f
C1040 VDPWR.n606 VGND 0.89889f
C1041 VDPWR.n607 VGND 1.33585f
C1042 VDPWR.n608 VGND 0.98231f
C1043 VDPWR.n609 VGND 0.04096f
C1044 VDPWR.n610 VGND 0.10703f
C1045 VDPWR.n611 VGND 0.11157f
C1046 VDPWR.n612 VGND 0.01923f
C1047 VDPWR.n613 VGND 0.35958f
C1048 VDPWR.n614 VGND 0.65864f
C1049 VDPWR.n615 VGND 0.20877f
C1050 VDPWR.n616 VGND 0.02935f
C1051 VDPWR.n617 VGND 0.03179f
C1052 VDPWR.n618 VGND 1.26615f
C1053 VDPWR.n619 VGND 1.09499f
C1054 VDPWR.n620 VGND 0.04105f
C1055 VDPWR.n621 VGND 0.04173f
C1056 VDPWR.n622 VGND 0.37096f
C1057 VDPWR.n623 VGND 0.0058f
C1058 VDPWR.n624 VGND 0.04097f
C1059 VDPWR.n625 VGND 0.20177f
C1060 VDPWR.n626 VGND 1.28429f
C1061 VDPWR.n627 VGND 0.03179f
C1062 VDPWR.n628 VGND 0.02931f
C1063 VDPWR.n629 VGND 0.01419f
C1064 VDPWR.n630 VGND 0.03137f
C1065 VDPWR.n631 VGND 0.42215f
C1066 VDPWR.n632 VGND 0.31975f
C1067 VDPWR.n633 VGND 0.27303f
C1068 VDPWR.n634 VGND 1.61926f
C1069 VDPWR.n635 VGND 1.15572f
C1070 VDPWR.n636 VGND 4.12112f
C1071 VDPWR.n637 VGND 3.522f
C1072 VDPWR.n638 VGND 10.2724f
C1073 VDPWR.n639 VGND 11.9627f
C1074 VDPWR.n640 VGND 11.3695f
C1075 VDPWR.n641 VGND 10.2909f
C1076 VDPWR.n642 VGND 1.06447f
C1077 VDPWR.n643 VGND 0.44351f
C1078 VDPWR.n644 VGND 0.17688f
C1079 VDPWR.n645 VGND 0.44015f
C1080 VDPWR.n646 VGND 3.25132f
C1081 VDPWR.n647 VGND 2.27269f
C1082 VDPWR.n648 VGND 4.69038f
C1083 VDPWR.n649 VGND 3.13272f
C1084 VDPWR.n650 VGND 3.154f
C1085 VDPWR.n651 VGND 1.99355f
C1086 VDPWR.n652 VGND 0.00232f
C1087 VDPWR.n653 VGND 0.1363f
C1088 VDPWR.n654 VGND 0.00234f
C1089 VDPWR.n655 VGND 0.01025f
C1090 VDPWR.n656 VGND 0.0152f
C1091 VDPWR.n657 VGND 0.00977f
C1092 VDPWR.n658 VGND 0.0152f
C1093 VDPWR.n659 VGND 0.22879f
C1094 VDPWR.n660 VGND 0.01011f
C1095 VDPWR.n661 VGND 0.0152f
C1096 VDPWR.n662 VGND 0.22879f
C1097 VDPWR.n663 VGND 0.01558f
C1098 VDPWR.n664 VGND 0.01558f
C1099 VDPWR.n665 VGND 0.01519f
C1100 VDPWR.n666 VGND 0.00544f
C1101 VDPWR.n667 VGND 0.00544f
C1102 VDPWR.n668 VGND 0.10818f
C1103 VDPWR.n669 VGND 0.00781f
C1104 VDPWR.n670 VGND 0.01558f
C1105 VDPWR.n671 VGND 0.01558f
C1106 VDPWR.n672 VGND 0.22879f
C1107 VDPWR.n673 VGND 0.01558f
C1108 VDPWR.n674 VGND 0.01558f
C1109 VDPWR.n675 VGND 0.00781f
C1110 VDPWR.n676 VGND 0.01558f
C1111 VDPWR.n677 VGND 0.01558f
C1112 VDPWR.n678 VGND 0.00781f
C1113 VDPWR.n679 VGND 0.0152f
C1114 VDPWR.n680 VGND 0.01519f
C1115 VDPWR.n681 VGND 0.0152f
C1116 VDPWR.n682 VGND 0.0152f
C1117 VDPWR.n683 VGND 0.18969f
C1118 VDPWR.n684 VGND 0.0152f
C1119 VDPWR.n685 VGND 0.0152f
C1120 VDPWR.n686 VGND 0.18969f
C1121 VDPWR.n687 VGND 0.0152f
C1122 VDPWR.n688 VGND 0.0152f
C1123 VDPWR.n689 VGND 0.01519f
C1124 VDPWR.n690 VGND 0.0152f
C1125 VDPWR.n691 VGND 0.19114f
C1126 VDPWR.n692 VGND 0.0152f
C1127 VDPWR.n693 VGND 0.01519f
C1128 VDPWR.n694 VGND 0.00544f
C1129 VDPWR.n695 VGND 0.02419f
C1130 VDPWR.n696 VGND 0.10818f
C1131 VDPWR.n697 VGND 0.02433f
C1132 VDPWR.n698 VGND 0.00544f
C1133 VDPWR.n699 VGND 0.00781f
C1134 VDPWR.n700 VGND 0.0152f
C1135 VDPWR.n701 VGND 0.0152f
C1136 VDPWR.n702 VGND 0.19114f
C1137 VDPWR.n703 VGND 0.19114f
C1138 VDPWR.n704 VGND 0.01011f
C1139 VDPWR.n705 VGND 0.01025f
C1140 VDPWR.n706 VGND 0.00977f
C1141 VDPWR.n707 VGND 0.00977f
C1142 VDPWR.n708 VGND 0.00977f
C1143 VDPWR.n709 VGND 0.22879f
C1144 VDPWR.n710 VGND 0.00464f
C1145 VDPWR.n711 VGND 0.00464f
C1146 VDPWR.n712 VGND 0.00977f
C1147 VDPWR.n713 VGND 0.00977f
C1148 VDPWR.n714 VGND 0.01011f
C1149 VDPWR.n715 VGND 0.00977f
C1150 VDPWR.n716 VGND 0.01025f
C1151 VDPWR.n717 VGND 0.01025f
C1152 VDPWR.n718 VGND 0.00975f
C1153 VDPWR.n719 VGND 0.01011f
C1154 VDPWR.n720 VGND 0.0152f
C1155 VDPWR.n721 VGND 0.0152f
C1156 VDPWR.n722 VGND 0.00977f
C1157 VDPWR.n723 VGND 0.00977f
C1158 VDPWR.n724 VGND 0.0152f
C1159 VDPWR.n725 VGND 0.0152f
C1160 VDPWR.n726 VGND 0.22879f
C1161 VDPWR.n727 VGND 0.01011f
C1162 VDPWR.n728 VGND 0.01011f
C1163 VDPWR.n729 VGND 0.01025f
C1164 VDPWR.n730 VGND 0.00234f
C1165 VDPWR.n731 VGND 0.00544f
C1166 VDPWR.n732 VGND 0.00781f
C1167 VDPWR.n733 VGND 0.01558f
C1168 VDPWR.n734 VGND 0.01558f
C1169 VDPWR.n735 VGND 0.22879f
C1170 VDPWR.n736 VGND 0.01558f
C1171 VDPWR.n737 VGND 0.01558f
C1172 VDPWR.n738 VGND 0.00781f
C1173 VDPWR.n739 VGND 0.22879f
C1174 VDPWR.n740 VGND 0.0152f
C1175 VDPWR.n741 VGND 0.01558f
C1176 VDPWR.n742 VGND 0.01558f
C1177 VDPWR.n743 VGND 0.00544f
C1178 VDPWR.n744 VGND 0.00781f
C1179 VDPWR.n745 VGND 0.01558f
C1180 VDPWR.n746 VGND 0.01558f
C1181 VDPWR.n747 VGND 0.01519f
C1182 VDPWR.n748 VGND 0.10818f
C1183 VDPWR.n749 VGND 0.03898f
C1184 VDPWR.n750 VGND 0.00544f
C1185 VDPWR.n751 VGND 0.00781f
C1186 VDPWR.n752 VGND 0.0152f
C1187 VDPWR.n753 VGND 0.0152f
C1188 VDPWR.n754 VGND 0.19114f
C1189 VDPWR.n755 VGND 0.0152f
C1190 VDPWR.n756 VGND 0.0152f
C1191 VDPWR.n757 VGND 0.01519f
C1192 VDPWR.n758 VGND 0.0152f
C1193 VDPWR.n759 VGND 0.18969f
C1194 VDPWR.n760 VGND 0.0152f
C1195 VDPWR.n761 VGND 0.0152f
C1196 VDPWR.n762 VGND 0.18969f
C1197 VDPWR.n763 VGND 0.0152f
C1198 VDPWR.n764 VGND 0.0152f
C1199 VDPWR.n765 VGND 0.01519f
C1200 VDPWR.n766 VGND 0.0152f
C1201 VDPWR.n767 VGND 0.22879f
C1202 VDPWR.n768 VGND 0.01011f
C1203 VDPWR.n769 VGND 0.01011f
C1204 VDPWR.n770 VGND 0.00977f
C1205 VDPWR.n771 VGND 0.00977f
C1206 VDPWR.n772 VGND 0.00977f
C1207 VDPWR.n773 VGND 0.00464f
C1208 VDPWR.n774 VGND 0.22879f
C1209 VDPWR.n775 VGND 0.00977f
C1210 VDPWR.n776 VGND 0.01025f
C1211 VDPWR.n777 VGND 0.00977f
C1212 VDPWR.n778 VGND 0.00977f
C1213 VDPWR.n779 VGND 0.00464f
C1214 VDPWR.n780 VGND 0.22879f
C1215 VDPWR.n781 VGND 0.22879f
C1216 VDPWR.n782 VGND 0.01025f
C1217 VDPWR.n783 VGND 0.01025f
C1218 VDPWR.n784 VGND 0.00977f
C1219 VDPWR.n785 VGND 0.01011f
C1220 VDPWR.n786 VGND 0.0152f
C1221 VDPWR.n787 VGND 0.0152f
C1222 VDPWR.n788 VGND 0.19114f
C1223 VDPWR.n789 VGND 0.19114f
C1224 VDPWR.n790 VGND 0.0152f
C1225 VDPWR.n791 VGND 0.01519f
C1226 VDPWR.n792 VGND 0.00544f
C1227 VDPWR.n793 VGND 0.02419f
C1228 VDPWR.n794 VGND 0.10818f
C1229 VDPWR.n795 VGND 0.08633f
C1230 VDPWR.n796 VGND 0.06836f
C1231 VDPWR.n797 VGND 0.00232f
C1232 VDPWR.n798 VGND 0.00975f
C1233 VDPWR.n799 VGND 0.01011f
C1234 VDPWR.n800 VGND 0.0152f
C1235 VDPWR.n801 VGND 0.0152f
C1236 VDPWR.n802 VGND 0.19114f
C1237 VDPWR.n803 VGND 0.19114f
C1238 VDPWR.n804 VGND 0.01011f
C1239 VDPWR.n805 VGND 0.01011f
C1240 VDPWR.n806 VGND 0.0152f
C1241 VDPWR.n807 VGND 0.00977f
C1242 VDPWR.n808 VGND 0.01025f
C1243 VDPWR.n809 VGND 0.01025f
C1244 VDPWR.n810 VGND 0.00977f
C1245 VDPWR.n811 VGND 0.01011f
C1246 VDPWR.n812 VGND 0.0152f
C1247 VDPWR.n813 VGND 0.01011f
C1248 VDPWR.n814 VGND 0.22879f
C1249 VDPWR.n815 VGND 0.01011f
C1250 VDPWR.n816 VGND 0.00977f
C1251 VDPWR.n817 VGND 0.01025f
C1252 VDPWR.n818 VGND 0.01025f
C1253 VDPWR.n819 VGND 0.00977f
C1254 VDPWR.n820 VGND 0.00234f
C1255 VDPWR.n821 VGND 0.00464f
C1256 VDPWR.n822 VGND 0.22879f
C1257 VDPWR.n823 VGND 0.00464f
C1258 VDPWR.n824 VGND 0.00977f
C1259 VDPWR.n825 VGND 0.01011f
C1260 VDPWR.n826 VGND 0.22879f
C1261 VDPWR.n827 VGND 0.01011f
C1262 VDPWR.n828 VGND 0.01011f
C1263 VDPWR.n829 VGND 0.00975f
C1264 VDPWR.n830 VGND 0.00232f
C1265 VDPWR.n831 VGND 0.06815f
C1266 VDPWR.n832 VGND 0.03649f
C1267 VDPWR.n833 VGND 0.36064f
C1268 VDPWR.n834 VGND 0.29729f
C1269 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A VGND 0.74657f
C1270 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G VGND 0.61957f
C1271 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin VGND 0.52606f
C1272 uo_out[2] VGND 3.26277f
C1273 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin VGND 0.52606f
C1274 uo_out[1] VGND 1.87298f
C1275 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin VGND 0.52752f
C1276 uo_out[0] VGND 1.64603f
C1277 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin VGND 0.52606f
C1278 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out VGND 1.20912f
C1279 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin VGND 0.52707f
C1280 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out VGND 1.2937f
C1281 VDPWR VGND 0.45143p
C1282 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin VGND 0.54717f
C1283 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out VGND 1.40293f
C1284 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin VGND 0.52756f
C1285 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 VGND 0.22293f
C1286 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin VGND 0.52606f
C1287 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out VGND 0.28552f
C1288 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin VGND 0.52645f
C1289 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out VGND 0.30478f
C1290 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin VGND 0.53627f
C1291 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out VGND 0.45287f
C1292 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/m1_n100_n100# VGND 0.10852f
C1293 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VGND 1.29945f
C1294 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in VGND 0.81081f
C1295 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G VGND 0.55523f
C1296 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VGND 3.05906f
C1297 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B VGND 0.42095f
C1298 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G VGND 0.55051f
C1299 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G VGND 0.5548f
C1300 ua[0] VGND 70.23664f
C1301 flashADC_3bit_0/comp_p_6/tail VGND 1.94675f
C1302 flashADC_3bit_0/comp_p_6/vbias_p VGND 14.26128f
C1303 uio_out[1] VGND 12.2039f
C1304 flashADC_3bit_0/comp_p_6/latch_right VGND 3.82409f
C1305 flashADC_3bit_0/comp_p_6/out_left VGND 3.36247f
C1306 flashADC_3bit_0/comp_p_6/latch_left VGND 3.98416f
C1307 flashADC_3bit_0/comp_p_5/tail VGND 1.09616f
C1308 uio_out[0] VGND 14.97629f
C1309 flashADC_3bit_0/comp_p_5/latch_right VGND 3.4916f
C1310 flashADC_3bit_0/comp_p_5/out_left VGND 2.14956f
C1311 flashADC_3bit_0/comp_p_5/latch_left VGND 3.68553f
C1312 flashADC_3bit_0/comp_p_4/tail VGND 1.09616f
C1313 uo_out[7] VGND 12.0344f
C1314 flashADC_3bit_0/comp_p_4/latch_right VGND 3.4916f
C1315 flashADC_3bit_0/comp_p_4/out_left VGND 3.01907f
C1316 flashADC_3bit_0/comp_p_4/latch_left VGND 3.68553f
C1317 flashADC_3bit_0/comp_p_3/tail VGND 1.46483f
C1318 uo_out[6] VGND 10.30018f
C1319 flashADC_3bit_0/comp_p_3/latch_right VGND 3.54536f
C1320 flashADC_3bit_0/comp_p_3/out_left VGND 3.74413f
C1321 flashADC_3bit_0/comp_p_3/latch_left VGND 10.64134f
C1322 flashADC_3bit_0/comp_p_2/tail VGND 1.42426f
C1323 uo_out[5] VGND 9.89908f
C1324 flashADC_3bit_0/comp_p_2/latch_right VGND 3.52097f
C1325 flashADC_3bit_0/comp_p_2/out_left VGND 3.30109f
C1326 flashADC_3bit_0/comp_p_2/latch_left VGND 3.70871f
C1327 flashADC_3bit_0/comp_p_0/tail VGND 1.18403f
C1328 uo_out[4] VGND 8.01901f
C1329 flashADC_3bit_0/comp_p_0/latch_right VGND 3.50563f
C1330 flashADC_3bit_0/comp_p_0/out_left VGND 2.37299f
C1331 flashADC_3bit_0/comp_p_0/latch_left VGND 9.17593f
C1332 flashADC_3bit_0/comp_p_1/tail VGND 1.19602f
C1333 uo_out[3] VGND 7.65664f
C1334 flashADC_3bit_0/comp_p_1/latch_right VGND 3.50878f
C1335 flashADC_3bit_0/comp_p_1/out_left VGND 3.65291f
C1336 flashADC_3bit_0/comp_p_1/latch_left VGND 3.70233f
C1337 flashADC_3bit_0/comp_p_0/vinn VGND 5.25373f
C1338 flashADC_3bit_0/comp_p_2/vinn VGND 4.2345f
C1339 flashADC_3bit_0/comp_p_3/vinn VGND 7.45335f
C1340 flashADC_3bit_0/comp_p_4/vinn VGND 3.89664f
C1341 flashADC_3bit_0/comp_p_5/vinn VGND 4.82118f
C1342 flashADC_3bit_0/comp_p_6/vinn VGND 7.68303f
C1343 flashADC_3bit_0/comp_p_1/vinn VGND 5.90892f
C1344 ua[1] VGND 26.36458f
C1345 flashADC_3bit_0/vbias_generation_0/bias_n VGND 2.08206f
C1346 flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 VGND 1.64553f
C1347 flashADC_3bit_0/vbias_generation_0/XR_bias_3/R2 VGND 1.48055f
C1348 flashADC_3bit_0/vbias_generation_0/XR_bias_2/R2 VGND 1.59499f
.ends

