magic
tech sky130A
timestamp 1762644791
<< nwell >>
rect -100 -610 148 617
<< pmoslvt >>
rect -50 -500 50 500
<< pdiff >>
rect -79 494 -50 500
rect -79 -494 -73 494
rect -56 -494 -50 494
rect -79 -500 -50 -494
rect 50 494 79 500
rect 50 -494 56 494
rect 73 -494 79 494
rect 50 -500 79 -494
<< pdiffc >>
rect -73 -494 -56 494
rect 56 -494 73 494
<< nsubdiff >>
rect 113 536 130 568
rect 113 -574 130 -550
<< nsubdiffcont >>
rect 113 -550 130 536
<< poly >>
rect -50 541 50 549
rect -50 524 -42 541
rect 42 524 50 541
rect -50 500 50 524
rect -50 -524 50 -500
rect -50 -541 -42 -524
rect 42 -541 50 -524
rect -50 -549 50 -541
<< polycont >>
rect -42 524 42 541
rect -42 -541 42 -524
<< locali >>
rect -50 524 -42 541
rect 42 524 50 541
rect 113 536 130 568
rect -73 494 -56 502
rect -73 -502 -56 -494
rect 56 494 73 502
rect 56 -502 73 -494
rect -50 -541 -42 -524
rect 42 -541 50 -524
rect 113 -574 130 -550
<< viali >>
rect -42 524 42 541
rect -73 -494 -56 494
rect 56 -494 73 494
rect -42 -541 42 -524
<< metal1 >>
rect -48 541 48 544
rect -48 524 -42 541
rect 42 524 48 541
rect -48 521 48 524
rect -76 494 -53 500
rect -76 -494 -73 494
rect -56 -494 -53 494
rect -76 -500 -53 -494
rect 53 494 76 500
rect 53 -494 56 494
rect 73 -494 76 494
rect 53 -500 76 -494
rect -48 -524 48 -521
rect -48 -541 -42 -524
rect 42 -541 48 -524
rect -48 -544 48 -541
<< labels >>
rlabel pdiffc -64 0 -64 0 0 D
port 2 nsew
rlabel pdiffc 64 0 64 0 0 S
port 3 nsew
rlabel polycont 0 533 0 533 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -121 -583 121 583
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
