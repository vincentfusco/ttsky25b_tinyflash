VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tinyflash
  CLASS BLOCK ;
  FOREIGN tt_um_tinyflash ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 97.950996 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 11.940 216.710 105.060 221.200 ;
        RECT 11.940 203.590 27.070 216.710 ;
      LAYER nwell ;
        RECT 27.070 203.590 79.600 216.710 ;
      LAYER pwell ;
        RECT 79.600 212.520 85.180 216.710 ;
      LAYER nwell ;
        RECT 85.180 212.520 104.140 216.710 ;
      LAYER pwell ;
        RECT 104.140 212.520 105.060 216.710 ;
        RECT 79.600 206.320 105.060 212.520 ;
        RECT 79.600 203.590 85.180 206.320 ;
        RECT 11.940 197.940 85.180 203.590 ;
      LAYER nwell ;
        RECT 85.180 197.940 104.140 206.320 ;
      LAYER pwell ;
        RECT 104.140 197.940 105.060 206.320 ;
        RECT 105.610 206.150 106.040 207.320 ;
        RECT 11.940 194.840 105.060 197.940 ;
        RECT 107.100 197.760 107.530 198.930 ;
        RECT 11.940 194.550 100.670 194.840 ;
        RECT 102.920 194.550 105.060 194.840 ;
        RECT 11.940 192.810 105.060 194.550 ;
        RECT 11.940 166.570 27.070 192.810 ;
      LAYER nwell ;
        RECT 27.070 166.570 79.600 192.810 ;
      LAYER pwell ;
        RECT 79.600 191.740 105.060 192.810 ;
        RECT 79.600 183.360 85.180 191.740 ;
      LAYER nwell ;
        RECT 85.180 183.360 104.140 191.740 ;
      LAYER pwell ;
        RECT 104.140 183.360 105.060 191.740 ;
        RECT 79.600 177.160 105.060 183.360 ;
        RECT 79.600 168.780 85.180 177.160 ;
      LAYER nwell ;
        RECT 85.180 168.780 104.140 177.160 ;
      LAYER pwell ;
        RECT 104.140 168.780 105.060 177.160 ;
        RECT 79.600 166.570 105.060 168.780 ;
        RECT 11.940 155.790 105.060 166.570 ;
        RECT 11.940 145.470 50.810 155.790 ;
        RECT 11.940 142.670 37.980 145.470 ;
      LAYER nwell ;
        RECT 37.980 144.430 50.810 145.470 ;
        RECT 37.980 142.990 50.800 144.430 ;
        RECT 53.990 142.670 79.600 155.790 ;
      LAYER pwell ;
        RECT 79.600 142.670 105.060 155.790 ;
        RECT 11.940 141.170 105.060 142.670 ;
      LAYER li1 ;
        RECT 85.380 216.530 87.080 216.570 ;
        RECT 87.480 216.530 89.180 216.570 ;
        RECT 100.130 216.530 101.830 216.570 ;
        RECT 102.230 216.530 103.930 216.570 ;
        RECT 27.240 216.360 52.500 216.530 ;
        RECT 27.240 214.100 30.310 216.360 ;
        RECT 31.025 215.790 39.065 215.960 ;
        RECT 30.640 214.730 30.810 215.730 ;
        RECT 39.280 214.730 39.450 215.730 ;
        RECT 31.025 214.500 39.065 214.670 ;
        RECT 39.790 214.100 39.960 216.360 ;
        RECT 40.685 215.790 48.725 215.960 ;
        RECT 40.300 214.730 40.470 215.730 ;
        RECT 48.940 214.730 49.110 215.730 ;
        RECT 40.685 214.500 48.725 214.670 ;
        RECT 49.450 214.110 52.500 216.360 ;
        RECT 45.720 214.100 52.500 214.110 ;
        RECT 27.240 213.490 52.500 214.100 ;
        RECT 12.130 213.300 23.230 213.320 ;
        RECT 12.120 213.110 23.310 213.300 ;
        RECT 12.120 206.440 12.290 213.110 ;
        RECT 12.770 206.920 14.930 212.650 ;
        RECT 20.500 206.920 22.660 212.650 ;
        RECT 23.140 206.440 23.310 213.110 ;
        RECT 12.120 206.270 23.310 206.440 ;
        RECT 12.120 199.580 12.290 206.270 ;
        RECT 12.770 200.060 14.930 205.790 ;
        RECT 20.500 200.060 22.660 205.790 ;
        RECT 23.140 199.580 23.310 206.270 ;
        RECT 27.240 211.230 34.240 213.490 ;
        RECT 35.045 213.090 44.925 213.490 ;
        RECT 34.965 212.920 45.005 213.090 ;
        RECT 34.580 211.860 34.750 212.860 ;
        RECT 45.220 211.860 45.390 212.860 ;
        RECT 34.965 211.630 45.005 211.800 ;
        RECT 45.720 211.230 52.500 213.490 ;
        RECT 27.240 210.150 52.500 211.230 ;
        RECT 27.240 205.080 28.600 210.150 ;
        RECT 29.175 209.650 39.210 209.820 ;
        RECT 28.790 209.240 28.960 209.590 ;
        RECT 39.425 209.240 39.595 209.590 ;
        RECT 29.175 209.010 39.210 209.180 ;
        RECT 29.175 208.450 39.210 208.620 ;
        RECT 28.790 208.040 28.960 208.390 ;
        RECT 39.425 208.040 39.595 208.390 ;
        RECT 29.175 207.810 39.210 207.980 ;
        RECT 29.175 207.250 39.210 207.420 ;
        RECT 28.790 206.840 28.960 207.190 ;
        RECT 39.425 206.840 39.595 207.190 ;
        RECT 29.175 206.610 39.210 206.780 ;
        RECT 29.175 206.050 39.210 206.220 ;
        RECT 28.790 205.640 28.960 205.990 ;
        RECT 39.425 205.640 39.595 205.990 ;
        RECT 29.175 205.410 39.210 205.580 ;
        RECT 39.790 205.080 39.960 210.150 ;
        RECT 40.535 209.650 50.570 209.820 ;
        RECT 40.150 209.240 40.320 209.590 ;
        RECT 49.810 209.180 50.530 209.260 ;
        RECT 50.785 209.240 50.955 209.590 ;
        RECT 40.535 209.010 50.570 209.180 ;
        RECT 49.810 208.920 50.530 209.010 ;
        RECT 40.535 208.450 50.570 208.620 ;
        RECT 40.150 208.040 40.320 208.390 ;
        RECT 50.785 208.040 50.955 208.390 ;
        RECT 40.535 207.810 50.570 207.980 ;
        RECT 40.535 207.250 50.570 207.420 ;
        RECT 40.150 206.840 40.320 207.190 ;
        RECT 49.810 206.780 50.530 206.860 ;
        RECT 50.785 206.840 50.955 207.190 ;
        RECT 40.535 206.610 50.570 206.780 ;
        RECT 49.810 206.520 50.530 206.610 ;
        RECT 40.535 206.050 50.570 206.220 ;
        RECT 40.150 205.640 40.320 205.990 ;
        RECT 50.785 205.640 50.955 205.990 ;
        RECT 40.535 205.410 50.570 205.580 ;
        RECT 51.145 205.080 52.500 210.150 ;
        RECT 27.240 204.910 52.500 205.080 ;
        RECT 54.160 216.360 79.420 216.530 ;
        RECT 54.160 214.100 57.230 216.360 ;
        RECT 57.945 215.790 65.985 215.960 ;
        RECT 57.560 214.730 57.730 215.730 ;
        RECT 66.200 214.730 66.370 215.730 ;
        RECT 57.945 214.500 65.985 214.670 ;
        RECT 66.710 214.100 66.880 216.360 ;
        RECT 67.605 215.790 75.645 215.960 ;
        RECT 67.220 214.730 67.390 215.730 ;
        RECT 75.860 214.730 76.030 215.730 ;
        RECT 67.605 214.500 75.645 214.670 ;
        RECT 76.370 214.110 79.420 216.360 ;
        RECT 72.640 214.100 79.420 214.110 ;
        RECT 54.160 213.490 79.420 214.100 ;
        RECT 54.160 211.230 61.160 213.490 ;
        RECT 61.965 213.090 71.845 213.490 ;
        RECT 61.885 212.920 71.925 213.090 ;
        RECT 61.500 211.860 61.670 212.860 ;
        RECT 72.140 211.860 72.310 212.860 ;
        RECT 61.885 211.630 71.925 211.800 ;
        RECT 72.640 211.230 79.420 213.490 ;
        RECT 85.360 216.360 87.110 216.530 ;
        RECT 85.360 212.870 85.530 216.360 ;
        RECT 86.070 215.850 86.400 216.020 ;
        RECT 85.930 213.595 86.100 215.635 ;
        RECT 86.370 213.595 86.540 215.635 ;
        RECT 86.070 213.210 86.400 213.380 ;
        RECT 86.940 212.870 87.110 216.360 ;
        RECT 85.360 212.700 87.110 212.870 ;
        RECT 87.460 216.360 89.210 216.530 ;
        RECT 87.460 212.870 87.630 216.360 ;
        RECT 88.170 215.850 88.500 216.020 ;
        RECT 88.030 213.595 88.200 215.635 ;
        RECT 88.470 213.595 88.640 215.635 ;
        RECT 88.170 213.210 88.500 213.380 ;
        RECT 89.040 212.870 89.210 216.360 ;
        RECT 87.460 212.700 89.210 212.870 ;
        RECT 89.570 216.360 94.480 216.530 ;
        RECT 89.570 212.870 89.740 216.360 ;
        RECT 90.280 215.850 90.610 216.020 ;
        RECT 90.140 213.595 90.310 215.635 ;
        RECT 90.580 213.595 90.750 215.635 ;
        RECT 90.280 213.210 90.610 213.380 ;
        RECT 91.150 212.870 91.320 216.360 ;
        RECT 91.860 215.850 92.190 216.020 ;
        RECT 91.720 213.595 91.890 215.635 ;
        RECT 92.160 213.595 92.330 215.635 ;
        RECT 91.860 213.210 92.190 213.380 ;
        RECT 92.730 212.870 92.900 216.360 ;
        RECT 93.440 215.850 93.770 216.020 ;
        RECT 93.300 213.595 93.470 215.635 ;
        RECT 93.740 213.595 93.910 215.635 ;
        RECT 93.440 213.210 93.770 213.380 ;
        RECT 94.310 212.870 94.480 216.360 ;
        RECT 89.570 212.700 94.480 212.870 ;
        RECT 100.110 216.360 101.860 216.530 ;
        RECT 100.110 212.870 100.280 216.360 ;
        RECT 100.820 215.850 101.150 216.020 ;
        RECT 100.680 213.595 100.850 215.635 ;
        RECT 101.120 213.595 101.290 215.635 ;
        RECT 100.820 213.210 101.150 213.380 ;
        RECT 101.690 212.870 101.860 216.360 ;
        RECT 100.110 212.700 101.860 212.870 ;
        RECT 102.210 216.360 103.960 216.530 ;
        RECT 102.210 212.870 102.380 216.360 ;
        RECT 102.920 215.850 103.250 216.020 ;
        RECT 102.780 213.595 102.950 215.635 ;
        RECT 103.220 213.595 103.390 215.635 ;
        RECT 102.920 213.210 103.250 213.380 ;
        RECT 103.790 212.870 103.960 216.360 ;
        RECT 102.210 212.700 103.960 212.870 ;
        RECT 54.160 210.150 79.420 211.230 ;
        RECT 54.160 205.080 55.520 210.150 ;
        RECT 56.095 209.650 66.130 209.820 ;
        RECT 55.710 209.240 55.880 209.590 ;
        RECT 66.345 209.240 66.515 209.590 ;
        RECT 56.095 209.010 66.130 209.180 ;
        RECT 56.095 208.450 66.130 208.620 ;
        RECT 55.710 208.040 55.880 208.390 ;
        RECT 66.345 208.040 66.515 208.390 ;
        RECT 56.095 207.810 66.130 207.980 ;
        RECT 56.095 207.250 66.130 207.420 ;
        RECT 55.710 206.840 55.880 207.190 ;
        RECT 66.345 206.840 66.515 207.190 ;
        RECT 56.095 206.610 66.130 206.780 ;
        RECT 56.095 206.050 66.130 206.220 ;
        RECT 55.710 205.640 55.880 205.990 ;
        RECT 66.345 205.640 66.515 205.990 ;
        RECT 56.095 205.410 66.130 205.580 ;
        RECT 66.710 205.080 66.880 210.150 ;
        RECT 67.455 209.650 77.490 209.820 ;
        RECT 67.070 209.240 67.240 209.590 ;
        RECT 76.730 209.180 77.450 209.260 ;
        RECT 77.705 209.240 77.875 209.590 ;
        RECT 67.455 209.010 77.490 209.180 ;
        RECT 76.730 208.920 77.450 209.010 ;
        RECT 67.455 208.450 77.490 208.620 ;
        RECT 67.070 208.040 67.240 208.390 ;
        RECT 77.705 208.040 77.875 208.390 ;
        RECT 67.455 207.810 77.490 207.980 ;
        RECT 67.455 207.250 77.490 207.420 ;
        RECT 67.070 206.840 67.240 207.190 ;
        RECT 76.730 206.780 77.450 206.860 ;
        RECT 77.705 206.840 77.875 207.190 ;
        RECT 67.455 206.610 77.490 206.780 ;
        RECT 76.730 206.520 77.450 206.610 ;
        RECT 67.455 206.050 77.490 206.220 ;
        RECT 67.070 205.640 67.240 205.990 ;
        RECT 77.705 205.640 77.875 205.990 ;
        RECT 67.455 205.410 77.490 205.580 ;
        RECT 78.065 205.080 79.420 210.150 ;
        RECT 85.360 212.170 87.110 212.340 ;
        RECT 85.360 209.770 85.530 212.170 ;
        RECT 86.070 211.660 86.400 211.830 ;
        RECT 85.930 210.450 86.100 211.490 ;
        RECT 86.370 210.450 86.540 211.490 ;
        RECT 86.070 210.110 86.400 210.280 ;
        RECT 86.940 209.770 87.110 212.170 ;
        RECT 85.360 209.600 87.110 209.770 ;
        RECT 87.460 212.170 89.210 212.340 ;
        RECT 87.460 209.770 87.630 212.170 ;
        RECT 88.170 211.660 88.500 211.830 ;
        RECT 88.030 210.450 88.200 211.490 ;
        RECT 88.470 210.450 88.640 211.490 ;
        RECT 88.170 210.110 88.500 210.280 ;
        RECT 89.040 209.770 89.210 212.170 ;
        RECT 87.460 209.600 89.210 209.770 ;
        RECT 89.570 212.170 94.480 212.340 ;
        RECT 89.570 209.770 89.740 212.170 ;
        RECT 90.280 211.660 90.610 211.830 ;
        RECT 90.140 210.450 90.310 211.490 ;
        RECT 90.580 210.450 90.750 211.490 ;
        RECT 90.280 210.110 90.610 210.280 ;
        RECT 91.150 209.770 91.320 212.170 ;
        RECT 91.860 211.660 92.190 211.830 ;
        RECT 91.720 210.450 91.890 211.490 ;
        RECT 92.160 210.450 92.330 211.490 ;
        RECT 91.860 210.110 92.190 210.280 ;
        RECT 92.730 209.770 92.900 212.170 ;
        RECT 93.440 211.660 93.770 211.830 ;
        RECT 93.300 210.450 93.470 211.490 ;
        RECT 93.740 210.450 93.910 211.490 ;
        RECT 93.440 210.110 93.770 210.280 ;
        RECT 94.310 209.770 94.480 212.170 ;
        RECT 89.570 209.690 94.480 209.770 ;
        RECT 100.110 212.170 101.860 212.340 ;
        RECT 100.110 209.770 100.280 212.170 ;
        RECT 100.820 211.660 101.150 211.830 ;
        RECT 100.680 210.450 100.850 211.490 ;
        RECT 101.120 210.450 101.290 211.490 ;
        RECT 100.820 210.110 101.150 210.280 ;
        RECT 101.690 209.770 101.860 212.170 ;
        RECT 89.570 209.600 94.490 209.690 ;
        RECT 100.110 209.600 101.860 209.770 ;
        RECT 102.210 212.170 103.960 212.340 ;
        RECT 102.210 209.770 102.380 212.170 ;
        RECT 102.920 211.660 103.250 211.830 ;
        RECT 102.780 210.450 102.950 211.490 ;
        RECT 103.220 210.450 103.390 211.490 ;
        RECT 102.920 210.110 103.250 210.280 ;
        RECT 103.790 209.770 103.960 212.170 ;
        RECT 102.210 209.600 103.960 209.770 ;
        RECT 85.380 209.570 87.080 209.600 ;
        RECT 87.480 209.570 89.180 209.600 ;
        RECT 89.650 209.520 94.490 209.600 ;
        RECT 100.130 209.570 101.830 209.600 ;
        RECT 102.230 209.570 103.930 209.600 ;
        RECT 85.380 209.240 87.080 209.270 ;
        RECT 87.480 209.240 89.180 209.270 ;
        RECT 89.650 209.240 94.490 209.320 ;
        RECT 94.920 209.240 99.760 209.320 ;
        RECT 100.130 209.240 101.830 209.270 ;
        RECT 102.230 209.240 103.930 209.270 ;
        RECT 85.360 209.070 87.110 209.240 ;
        RECT 85.360 206.670 85.530 209.070 ;
        RECT 86.070 208.560 86.400 208.730 ;
        RECT 85.930 207.350 86.100 208.390 ;
        RECT 86.370 207.350 86.540 208.390 ;
        RECT 86.070 207.010 86.400 207.180 ;
        RECT 86.940 206.670 87.110 209.070 ;
        RECT 85.360 206.500 87.110 206.670 ;
        RECT 87.460 209.070 89.210 209.240 ;
        RECT 87.460 206.670 87.630 209.070 ;
        RECT 88.170 208.560 88.500 208.730 ;
        RECT 88.030 207.350 88.200 208.390 ;
        RECT 88.470 207.350 88.640 208.390 ;
        RECT 88.170 207.010 88.500 207.180 ;
        RECT 89.040 206.670 89.210 209.070 ;
        RECT 87.460 206.500 89.210 206.670 ;
        RECT 89.570 209.150 94.490 209.240 ;
        RECT 94.840 209.150 99.760 209.240 ;
        RECT 89.570 209.070 94.480 209.150 ;
        RECT 89.570 206.670 89.740 209.070 ;
        RECT 90.280 208.560 90.610 208.730 ;
        RECT 90.140 207.350 90.310 208.390 ;
        RECT 90.580 207.350 90.750 208.390 ;
        RECT 90.280 207.010 90.610 207.180 ;
        RECT 91.150 206.670 91.320 209.070 ;
        RECT 91.860 208.560 92.190 208.730 ;
        RECT 91.720 207.350 91.890 208.390 ;
        RECT 92.160 207.350 92.330 208.390 ;
        RECT 91.860 207.010 92.190 207.180 ;
        RECT 92.730 206.670 92.900 209.070 ;
        RECT 93.440 208.560 93.770 208.730 ;
        RECT 93.300 207.350 93.470 208.390 ;
        RECT 93.740 207.350 93.910 208.390 ;
        RECT 93.440 207.010 93.770 207.180 ;
        RECT 94.310 206.670 94.480 209.070 ;
        RECT 89.570 206.500 94.480 206.670 ;
        RECT 94.840 209.070 99.750 209.150 ;
        RECT 94.840 206.670 95.010 209.070 ;
        RECT 95.550 208.560 95.880 208.730 ;
        RECT 95.410 207.350 95.580 208.390 ;
        RECT 95.850 207.350 96.020 208.390 ;
        RECT 95.550 207.010 95.880 207.180 ;
        RECT 96.420 206.670 96.590 209.070 ;
        RECT 97.130 208.560 97.460 208.730 ;
        RECT 96.990 207.350 97.160 208.390 ;
        RECT 97.430 207.350 97.600 208.390 ;
        RECT 97.130 207.010 97.460 207.180 ;
        RECT 98.000 206.670 98.170 209.070 ;
        RECT 98.710 208.560 99.040 208.730 ;
        RECT 98.570 207.350 98.740 208.390 ;
        RECT 99.010 207.350 99.180 208.390 ;
        RECT 98.710 207.010 99.040 207.180 ;
        RECT 99.580 206.670 99.750 209.070 ;
        RECT 94.840 206.500 99.750 206.670 ;
        RECT 100.110 209.070 101.860 209.240 ;
        RECT 100.110 206.670 100.280 209.070 ;
        RECT 100.820 208.560 101.150 208.730 ;
        RECT 100.680 207.350 100.850 208.390 ;
        RECT 101.120 207.350 101.290 208.390 ;
        RECT 100.820 207.010 101.150 207.180 ;
        RECT 101.690 206.670 101.860 209.070 ;
        RECT 100.110 206.500 101.860 206.670 ;
        RECT 102.210 209.070 103.960 209.240 ;
        RECT 102.210 206.670 102.380 209.070 ;
        RECT 102.920 208.560 103.250 208.730 ;
        RECT 102.780 207.350 102.950 208.390 ;
        RECT 103.220 207.350 103.390 208.390 ;
        RECT 102.920 207.010 103.250 207.180 ;
        RECT 103.790 206.670 103.960 209.070 ;
        RECT 102.210 206.500 103.960 206.670 ;
        RECT 54.160 204.910 79.420 205.080 ;
        RECT 85.360 205.970 87.110 206.140 ;
        RECT 27.250 203.240 52.500 203.410 ;
        RECT 27.250 201.390 27.420 203.240 ;
        RECT 28.100 202.670 32.140 202.840 ;
        RECT 27.760 201.610 27.930 202.610 ;
        RECT 32.310 201.610 32.480 202.610 ;
        RECT 28.180 201.550 32.060 201.580 ;
        RECT 28.100 201.390 32.140 201.550 ;
        RECT 32.820 201.390 32.990 203.240 ;
        RECT 33.950 202.670 38.990 202.840 ;
        RECT 33.610 201.610 33.780 202.610 ;
        RECT 39.160 201.610 39.330 202.610 ;
        RECT 33.950 201.390 38.990 201.550 ;
        RECT 39.790 201.390 39.960 203.240 ;
        RECT 40.920 202.670 45.960 202.840 ;
        RECT 40.580 201.610 40.750 202.610 ;
        RECT 46.130 201.610 46.300 202.610 ;
        RECT 40.920 201.390 45.960 201.550 ;
        RECT 46.760 201.390 46.930 203.240 ;
        RECT 47.610 202.670 51.650 202.840 ;
        RECT 47.270 201.610 47.440 202.610 ;
        RECT 51.820 201.610 51.990 202.610 ;
        RECT 47.690 201.550 51.570 201.580 ;
        RECT 47.610 201.390 51.650 201.550 ;
        RECT 52.330 201.390 52.500 203.240 ;
        RECT 54.170 203.240 79.420 203.410 ;
        RECT 54.170 201.390 54.340 203.240 ;
        RECT 55.020 202.670 59.060 202.840 ;
        RECT 54.680 201.610 54.850 202.610 ;
        RECT 59.230 201.610 59.400 202.610 ;
        RECT 55.100 201.550 58.980 201.580 ;
        RECT 55.020 201.390 59.060 201.550 ;
        RECT 59.740 201.390 59.910 203.240 ;
        RECT 60.870 202.670 65.910 202.840 ;
        RECT 60.530 201.610 60.700 202.610 ;
        RECT 66.080 201.610 66.250 202.610 ;
        RECT 60.870 201.390 65.910 201.550 ;
        RECT 66.710 201.390 66.880 203.240 ;
        RECT 67.840 202.670 72.880 202.840 ;
        RECT 67.500 201.610 67.670 202.610 ;
        RECT 73.050 201.610 73.220 202.610 ;
        RECT 67.840 201.390 72.880 201.550 ;
        RECT 73.680 201.390 73.850 203.240 ;
        RECT 74.530 202.670 78.570 202.840 ;
        RECT 74.190 201.610 74.360 202.610 ;
        RECT 78.740 201.610 78.910 202.610 ;
        RECT 74.610 201.550 78.490 201.580 ;
        RECT 74.530 201.390 78.570 201.550 ;
        RECT 79.250 201.390 79.420 203.240 ;
        RECT 85.360 202.480 85.530 205.970 ;
        RECT 86.070 205.460 86.400 205.630 ;
        RECT 85.930 203.205 86.100 205.245 ;
        RECT 86.370 203.205 86.540 205.245 ;
        RECT 86.070 202.820 86.400 202.990 ;
        RECT 86.940 202.480 87.110 205.970 ;
        RECT 85.360 202.310 87.110 202.480 ;
        RECT 87.460 205.970 89.210 206.140 ;
        RECT 87.460 202.480 87.630 205.970 ;
        RECT 88.170 205.460 88.500 205.630 ;
        RECT 88.030 203.205 88.200 205.245 ;
        RECT 88.470 203.205 88.640 205.245 ;
        RECT 88.170 202.820 88.500 202.990 ;
        RECT 89.040 202.480 89.210 205.970 ;
        RECT 87.460 202.310 89.210 202.480 ;
        RECT 89.570 205.970 94.480 206.140 ;
        RECT 89.570 202.480 89.740 205.970 ;
        RECT 90.280 205.460 90.610 205.630 ;
        RECT 90.140 203.205 90.310 205.245 ;
        RECT 90.580 203.205 90.750 205.245 ;
        RECT 90.280 202.820 90.610 202.990 ;
        RECT 91.150 202.480 91.320 205.970 ;
        RECT 91.860 205.460 92.190 205.630 ;
        RECT 91.720 203.205 91.890 205.245 ;
        RECT 92.160 203.205 92.330 205.245 ;
        RECT 91.860 202.820 92.190 202.990 ;
        RECT 92.730 202.480 92.900 205.970 ;
        RECT 93.440 205.460 93.770 205.630 ;
        RECT 93.300 203.205 93.470 205.245 ;
        RECT 93.740 203.205 93.910 205.245 ;
        RECT 93.440 202.820 93.770 202.990 ;
        RECT 94.310 202.480 94.480 205.970 ;
        RECT 89.570 202.310 94.480 202.480 ;
        RECT 94.840 205.970 99.750 206.140 ;
        RECT 94.840 202.480 95.010 205.970 ;
        RECT 95.550 205.460 95.880 205.630 ;
        RECT 95.410 203.205 95.580 205.245 ;
        RECT 95.850 203.205 96.020 205.245 ;
        RECT 95.550 202.820 95.880 202.990 ;
        RECT 96.420 202.480 96.590 205.970 ;
        RECT 97.130 205.460 97.460 205.630 ;
        RECT 96.990 203.205 97.160 205.245 ;
        RECT 97.430 203.205 97.600 205.245 ;
        RECT 97.130 202.820 97.460 202.990 ;
        RECT 98.000 202.480 98.170 205.970 ;
        RECT 98.710 205.460 99.040 205.630 ;
        RECT 98.570 203.205 98.740 205.245 ;
        RECT 99.010 203.205 99.180 205.245 ;
        RECT 98.710 202.820 99.040 202.990 ;
        RECT 99.580 202.480 99.750 205.970 ;
        RECT 94.840 202.310 99.750 202.480 ;
        RECT 100.110 205.970 101.860 206.140 ;
        RECT 100.110 202.480 100.280 205.970 ;
        RECT 100.820 205.460 101.150 205.630 ;
        RECT 100.680 203.205 100.850 205.245 ;
        RECT 101.120 203.205 101.290 205.245 ;
        RECT 100.820 202.820 101.150 202.990 ;
        RECT 101.690 202.480 101.860 205.970 ;
        RECT 100.110 202.310 101.860 202.480 ;
        RECT 102.210 205.970 103.960 206.140 ;
        RECT 102.210 202.480 102.380 205.970 ;
        RECT 102.920 205.460 103.250 205.630 ;
        RECT 102.780 203.205 102.950 205.245 ;
        RECT 103.220 203.205 103.390 205.245 ;
        RECT 102.920 202.820 103.250 202.990 ;
        RECT 103.790 202.480 103.960 205.970 ;
        RECT 102.210 202.310 103.960 202.480 ;
        RECT 85.380 202.270 87.080 202.310 ;
        RECT 87.480 202.270 89.180 202.310 ;
        RECT 100.130 202.270 101.830 202.310 ;
        RECT 102.230 202.270 103.930 202.310 ;
        RECT 85.380 201.950 87.080 201.990 ;
        RECT 87.480 201.950 89.180 201.990 ;
        RECT 100.130 201.950 101.830 201.990 ;
        RECT 102.230 201.950 103.930 201.990 ;
        RECT 12.120 199.410 23.310 199.580 ;
        RECT 12.120 192.720 12.290 199.410 ;
        RECT 12.770 193.200 14.930 198.930 ;
        RECT 20.500 193.200 22.660 198.930 ;
        RECT 23.140 192.720 23.310 199.410 ;
        RECT 27.240 200.810 52.500 201.390 ;
        RECT 27.240 198.550 32.990 200.810 ;
        RECT 33.950 200.240 38.990 200.410 ;
        RECT 33.610 199.180 33.780 200.180 ;
        RECT 39.160 199.180 39.330 200.180 ;
        RECT 33.950 198.950 38.990 199.120 ;
        RECT 39.790 198.550 39.960 200.810 ;
        RECT 40.920 200.240 45.960 200.410 ;
        RECT 40.580 199.180 40.750 200.180 ;
        RECT 46.130 199.180 46.300 200.180 ;
        RECT 40.920 198.950 45.960 199.120 ;
        RECT 46.760 198.550 52.500 200.810 ;
        RECT 27.240 198.380 52.500 198.550 ;
        RECT 54.160 200.810 79.420 201.390 ;
        RECT 54.160 198.550 59.910 200.810 ;
        RECT 60.870 200.240 65.910 200.410 ;
        RECT 60.530 199.180 60.700 200.180 ;
        RECT 66.080 199.180 66.250 200.180 ;
        RECT 60.870 198.950 65.910 199.120 ;
        RECT 66.710 198.550 66.880 200.810 ;
        RECT 67.840 200.240 72.880 200.410 ;
        RECT 67.500 199.180 67.670 200.180 ;
        RECT 73.050 199.180 73.220 200.180 ;
        RECT 67.840 198.950 72.880 199.120 ;
        RECT 73.680 198.550 79.420 200.810 ;
        RECT 54.160 198.380 79.420 198.550 ;
        RECT 85.360 201.780 87.110 201.950 ;
        RECT 85.360 198.290 85.530 201.780 ;
        RECT 86.070 201.270 86.400 201.440 ;
        RECT 85.930 199.015 86.100 201.055 ;
        RECT 86.370 199.015 86.540 201.055 ;
        RECT 86.070 198.630 86.400 198.800 ;
        RECT 86.940 198.290 87.110 201.780 ;
        RECT 85.360 198.120 87.110 198.290 ;
        RECT 87.460 201.780 89.210 201.950 ;
        RECT 87.460 198.290 87.630 201.780 ;
        RECT 88.170 201.270 88.500 201.440 ;
        RECT 88.030 199.015 88.200 201.055 ;
        RECT 88.470 199.015 88.640 201.055 ;
        RECT 88.170 198.630 88.500 198.800 ;
        RECT 89.040 198.290 89.210 201.780 ;
        RECT 87.460 198.120 89.210 198.290 ;
        RECT 89.570 201.780 94.480 201.950 ;
        RECT 89.570 198.290 89.740 201.780 ;
        RECT 90.280 201.270 90.610 201.440 ;
        RECT 90.140 199.015 90.310 201.055 ;
        RECT 90.580 199.015 90.750 201.055 ;
        RECT 90.280 198.630 90.610 198.800 ;
        RECT 91.150 198.290 91.320 201.780 ;
        RECT 91.860 201.270 92.190 201.440 ;
        RECT 91.720 199.015 91.890 201.055 ;
        RECT 92.160 199.015 92.330 201.055 ;
        RECT 91.860 198.630 92.190 198.800 ;
        RECT 92.730 198.290 92.900 201.780 ;
        RECT 93.440 201.270 93.770 201.440 ;
        RECT 93.300 199.015 93.470 201.055 ;
        RECT 93.740 199.015 93.910 201.055 ;
        RECT 93.440 198.630 93.770 198.800 ;
        RECT 94.310 198.290 94.480 201.780 ;
        RECT 89.570 198.120 94.480 198.290 ;
        RECT 100.110 201.780 101.860 201.950 ;
        RECT 100.110 198.290 100.280 201.780 ;
        RECT 100.820 201.270 101.150 201.440 ;
        RECT 100.680 199.015 100.850 201.055 ;
        RECT 101.120 199.015 101.290 201.055 ;
        RECT 100.820 198.630 101.150 198.800 ;
        RECT 101.690 198.290 101.860 201.780 ;
        RECT 100.110 198.120 101.860 198.290 ;
        RECT 102.210 201.780 103.960 201.950 ;
        RECT 102.210 198.290 102.380 201.780 ;
        RECT 102.920 201.270 103.250 201.440 ;
        RECT 102.780 199.015 102.950 201.055 ;
        RECT 103.220 199.015 103.390 201.055 ;
        RECT 102.920 198.630 103.250 198.800 ;
        RECT 103.790 198.290 103.960 201.780 ;
        RECT 102.210 198.120 103.960 198.290 ;
        RECT 27.240 197.850 52.500 198.020 ;
        RECT 27.240 195.590 32.990 197.850 ;
        RECT 33.950 197.280 38.990 197.450 ;
        RECT 33.610 196.220 33.780 197.220 ;
        RECT 39.160 196.220 39.330 197.220 ;
        RECT 33.950 195.990 38.990 196.160 ;
        RECT 39.790 195.590 39.960 197.850 ;
        RECT 40.920 197.280 45.960 197.450 ;
        RECT 40.580 196.220 40.750 197.220 ;
        RECT 46.130 196.220 46.300 197.220 ;
        RECT 40.920 195.990 45.960 196.160 ;
        RECT 46.760 195.590 52.500 197.850 ;
        RECT 27.240 195.010 52.500 195.590 ;
        RECT 54.160 197.850 79.420 198.020 ;
        RECT 54.160 195.590 59.910 197.850 ;
        RECT 60.870 197.280 65.910 197.450 ;
        RECT 60.530 196.220 60.700 197.220 ;
        RECT 66.080 196.220 66.250 197.220 ;
        RECT 60.870 195.990 65.910 196.160 ;
        RECT 66.710 195.590 66.880 197.850 ;
        RECT 67.840 197.280 72.880 197.450 ;
        RECT 67.500 196.220 67.670 197.220 ;
        RECT 73.050 196.220 73.220 197.220 ;
        RECT 67.840 195.990 72.880 196.160 ;
        RECT 73.680 195.590 79.420 197.850 ;
        RECT 54.160 195.010 79.420 195.590 ;
        RECT 85.360 197.590 87.110 197.760 ;
        RECT 85.360 195.190 85.530 197.590 ;
        RECT 86.070 197.080 86.400 197.250 ;
        RECT 85.930 195.870 86.100 196.910 ;
        RECT 86.370 195.870 86.540 196.910 ;
        RECT 86.070 195.530 86.400 195.700 ;
        RECT 86.940 195.190 87.110 197.590 ;
        RECT 85.360 195.020 87.110 195.190 ;
        RECT 87.460 197.590 89.210 197.760 ;
        RECT 87.460 195.190 87.630 197.590 ;
        RECT 88.170 197.080 88.500 197.250 ;
        RECT 88.030 195.870 88.200 196.910 ;
        RECT 88.470 195.870 88.640 196.910 ;
        RECT 88.170 195.530 88.500 195.700 ;
        RECT 89.040 195.190 89.210 197.590 ;
        RECT 87.460 195.020 89.210 195.190 ;
        RECT 89.570 197.590 94.480 197.760 ;
        RECT 89.570 195.190 89.740 197.590 ;
        RECT 90.280 197.080 90.610 197.250 ;
        RECT 90.140 195.870 90.310 196.910 ;
        RECT 90.580 195.870 90.750 196.910 ;
        RECT 90.280 195.530 90.610 195.700 ;
        RECT 91.150 195.190 91.320 197.590 ;
        RECT 91.860 197.080 92.190 197.250 ;
        RECT 91.720 195.870 91.890 196.910 ;
        RECT 92.160 195.870 92.330 196.910 ;
        RECT 91.860 195.530 92.190 195.700 ;
        RECT 92.730 195.190 92.900 197.590 ;
        RECT 93.440 197.080 93.770 197.250 ;
        RECT 93.300 195.870 93.470 196.910 ;
        RECT 93.740 195.870 93.910 196.910 ;
        RECT 93.440 195.530 93.770 195.700 ;
        RECT 94.310 195.190 94.480 197.590 ;
        RECT 89.570 195.110 94.480 195.190 ;
        RECT 100.110 197.590 101.860 197.760 ;
        RECT 100.110 195.190 100.280 197.590 ;
        RECT 100.820 197.080 101.150 197.250 ;
        RECT 100.680 195.870 100.850 196.910 ;
        RECT 101.120 195.870 101.290 196.910 ;
        RECT 100.820 195.530 101.150 195.700 ;
        RECT 101.690 195.190 101.860 197.590 ;
        RECT 89.570 195.020 94.490 195.110 ;
        RECT 100.110 195.020 101.860 195.190 ;
        RECT 102.210 197.590 103.960 197.760 ;
        RECT 102.210 195.190 102.380 197.590 ;
        RECT 102.920 197.080 103.250 197.250 ;
        RECT 102.780 195.870 102.950 196.910 ;
        RECT 103.220 195.870 103.390 196.910 ;
        RECT 102.920 195.530 103.250 195.700 ;
        RECT 103.790 195.190 103.960 197.590 ;
        RECT 102.210 195.020 103.960 195.190 ;
        RECT 27.250 193.160 27.420 195.010 ;
        RECT 28.100 194.850 32.140 195.010 ;
        RECT 28.180 194.820 32.060 194.850 ;
        RECT 27.760 193.790 27.930 194.790 ;
        RECT 32.310 193.790 32.480 194.790 ;
        RECT 28.100 193.560 32.140 193.730 ;
        RECT 32.820 193.160 32.990 195.010 ;
        RECT 33.950 194.850 38.990 195.010 ;
        RECT 33.610 193.790 33.780 194.790 ;
        RECT 39.160 193.790 39.330 194.790 ;
        RECT 33.950 193.560 38.990 193.730 ;
        RECT 39.790 193.160 39.960 195.010 ;
        RECT 40.920 194.850 45.960 195.010 ;
        RECT 40.580 193.790 40.750 194.790 ;
        RECT 46.130 193.790 46.300 194.790 ;
        RECT 40.920 193.560 45.960 193.730 ;
        RECT 46.760 193.160 46.930 195.010 ;
        RECT 47.610 194.850 51.650 195.010 ;
        RECT 47.690 194.820 51.570 194.850 ;
        RECT 47.270 193.790 47.440 194.790 ;
        RECT 51.820 193.790 51.990 194.790 ;
        RECT 47.610 193.560 51.650 193.730 ;
        RECT 52.330 193.160 52.500 195.010 ;
        RECT 27.250 192.990 52.500 193.160 ;
        RECT 54.170 193.160 54.340 195.010 ;
        RECT 55.020 194.850 59.060 195.010 ;
        RECT 55.100 194.820 58.980 194.850 ;
        RECT 54.680 193.790 54.850 194.790 ;
        RECT 59.230 193.790 59.400 194.790 ;
        RECT 55.020 193.560 59.060 193.730 ;
        RECT 59.740 193.160 59.910 195.010 ;
        RECT 60.870 194.850 65.910 195.010 ;
        RECT 60.530 193.790 60.700 194.790 ;
        RECT 66.080 193.790 66.250 194.790 ;
        RECT 60.870 193.560 65.910 193.730 ;
        RECT 66.710 193.160 66.880 195.010 ;
        RECT 67.840 194.850 72.880 195.010 ;
        RECT 67.500 193.790 67.670 194.790 ;
        RECT 73.050 193.790 73.220 194.790 ;
        RECT 67.840 193.560 72.880 193.730 ;
        RECT 73.680 193.160 73.850 195.010 ;
        RECT 74.530 194.850 78.570 195.010 ;
        RECT 74.610 194.820 78.490 194.850 ;
        RECT 74.190 193.790 74.360 194.790 ;
        RECT 78.740 193.790 78.910 194.790 ;
        RECT 74.530 193.560 78.570 193.730 ;
        RECT 79.250 193.160 79.420 195.010 ;
        RECT 85.380 194.990 87.080 195.020 ;
        RECT 87.480 194.990 89.180 195.020 ;
        RECT 89.650 194.940 94.490 195.020 ;
        RECT 100.130 194.990 101.830 195.020 ;
        RECT 102.230 194.990 103.930 195.020 ;
        RECT 85.380 194.660 87.080 194.690 ;
        RECT 87.480 194.660 89.180 194.690 ;
        RECT 54.170 192.990 79.420 193.160 ;
        RECT 85.360 194.490 87.110 194.660 ;
        RECT 12.120 192.550 23.310 192.720 ;
        RECT 12.120 185.860 12.290 192.550 ;
        RECT 12.770 186.340 14.930 192.070 ;
        RECT 20.500 186.340 22.660 192.070 ;
        RECT 23.140 185.860 23.310 192.550 ;
        RECT 85.360 192.090 85.530 194.490 ;
        RECT 86.070 193.980 86.400 194.150 ;
        RECT 85.930 192.770 86.100 193.810 ;
        RECT 86.370 192.770 86.540 193.810 ;
        RECT 86.070 192.430 86.400 192.600 ;
        RECT 86.940 192.090 87.110 194.490 ;
        RECT 85.360 191.920 87.110 192.090 ;
        RECT 87.460 194.490 89.210 194.660 ;
        RECT 87.460 192.090 87.630 194.490 ;
        RECT 88.170 193.980 88.500 194.150 ;
        RECT 88.030 192.770 88.200 193.810 ;
        RECT 88.470 192.770 88.640 193.810 ;
        RECT 88.170 192.430 88.500 192.600 ;
        RECT 89.040 192.090 89.210 194.490 ;
        RECT 87.460 191.920 89.210 192.090 ;
        RECT 12.120 185.690 23.310 185.860 ;
        RECT 12.120 179.000 12.290 185.690 ;
        RECT 12.770 179.480 14.930 185.210 ;
        RECT 20.500 179.480 22.660 185.210 ;
        RECT 23.140 179.000 23.310 185.690 ;
        RECT 27.240 191.320 52.500 191.490 ;
        RECT 27.240 186.250 28.600 191.320 ;
        RECT 29.175 190.820 39.210 190.990 ;
        RECT 28.790 190.410 28.960 190.760 ;
        RECT 39.425 190.410 39.595 190.760 ;
        RECT 29.175 190.180 39.210 190.350 ;
        RECT 29.175 189.620 39.210 189.790 ;
        RECT 28.790 189.210 28.960 189.560 ;
        RECT 39.425 189.210 39.595 189.560 ;
        RECT 29.175 188.980 39.210 189.150 ;
        RECT 29.175 188.420 39.210 188.590 ;
        RECT 28.790 188.010 28.960 188.360 ;
        RECT 39.425 188.010 39.595 188.360 ;
        RECT 29.175 187.780 39.210 187.950 ;
        RECT 29.175 187.220 39.210 187.390 ;
        RECT 28.790 186.810 28.960 187.160 ;
        RECT 39.425 186.810 39.595 187.160 ;
        RECT 29.175 186.580 39.210 186.750 ;
        RECT 39.790 186.250 39.960 191.320 ;
        RECT 40.535 190.820 50.570 190.990 ;
        RECT 40.150 190.410 40.320 190.760 ;
        RECT 50.785 190.410 50.955 190.760 ;
        RECT 40.535 190.180 50.570 190.350 ;
        RECT 49.810 189.790 50.530 189.880 ;
        RECT 40.535 189.620 50.570 189.790 ;
        RECT 40.150 189.210 40.320 189.560 ;
        RECT 49.810 189.540 50.530 189.620 ;
        RECT 50.785 189.210 50.955 189.560 ;
        RECT 40.535 188.980 50.570 189.150 ;
        RECT 40.535 188.420 50.570 188.590 ;
        RECT 40.150 188.010 40.320 188.360 ;
        RECT 50.785 188.010 50.955 188.360 ;
        RECT 40.535 187.780 50.570 187.950 ;
        RECT 49.810 187.390 50.530 187.480 ;
        RECT 40.535 187.220 50.570 187.390 ;
        RECT 40.150 186.810 40.320 187.160 ;
        RECT 49.810 187.140 50.530 187.220 ;
        RECT 50.785 186.810 50.955 187.160 ;
        RECT 40.535 186.580 50.570 186.750 ;
        RECT 51.145 186.250 52.500 191.320 ;
        RECT 27.240 185.170 52.500 186.250 ;
        RECT 27.240 182.910 34.240 185.170 ;
        RECT 34.965 184.600 45.005 184.770 ;
        RECT 34.580 183.540 34.750 184.540 ;
        RECT 45.220 183.540 45.390 184.540 ;
        RECT 34.965 183.310 45.005 183.480 ;
        RECT 35.045 182.910 44.925 183.310 ;
        RECT 45.720 182.910 52.500 185.170 ;
        RECT 27.240 182.300 52.500 182.910 ;
        RECT 27.240 180.040 30.310 182.300 ;
        RECT 31.025 181.730 39.065 181.900 ;
        RECT 30.640 180.670 30.810 181.670 ;
        RECT 39.280 180.670 39.450 181.670 ;
        RECT 31.025 180.440 39.065 180.610 ;
        RECT 39.790 180.040 39.960 182.300 ;
        RECT 45.720 182.290 52.500 182.300 ;
        RECT 40.685 181.730 48.725 181.900 ;
        RECT 40.300 180.670 40.470 181.670 ;
        RECT 48.940 180.670 49.110 181.670 ;
        RECT 40.685 180.440 48.725 180.610 ;
        RECT 49.450 180.040 52.500 182.290 ;
        RECT 27.240 179.870 52.500 180.040 ;
        RECT 54.160 191.320 79.420 191.490 ;
        RECT 54.160 186.250 55.520 191.320 ;
        RECT 56.095 190.820 66.130 190.990 ;
        RECT 55.710 190.410 55.880 190.760 ;
        RECT 66.345 190.410 66.515 190.760 ;
        RECT 56.095 190.180 66.130 190.350 ;
        RECT 56.095 189.620 66.130 189.790 ;
        RECT 55.710 189.210 55.880 189.560 ;
        RECT 66.345 189.210 66.515 189.560 ;
        RECT 56.095 188.980 66.130 189.150 ;
        RECT 56.095 188.420 66.130 188.590 ;
        RECT 55.710 188.010 55.880 188.360 ;
        RECT 66.345 188.010 66.515 188.360 ;
        RECT 56.095 187.780 66.130 187.950 ;
        RECT 56.095 187.220 66.130 187.390 ;
        RECT 55.710 186.810 55.880 187.160 ;
        RECT 66.345 186.810 66.515 187.160 ;
        RECT 56.095 186.580 66.130 186.750 ;
        RECT 66.710 186.250 66.880 191.320 ;
        RECT 67.455 190.820 77.490 190.990 ;
        RECT 67.070 190.410 67.240 190.760 ;
        RECT 77.705 190.410 77.875 190.760 ;
        RECT 67.455 190.180 77.490 190.350 ;
        RECT 76.730 189.790 77.450 189.880 ;
        RECT 67.455 189.620 77.490 189.790 ;
        RECT 67.070 189.210 67.240 189.560 ;
        RECT 76.730 189.540 77.450 189.620 ;
        RECT 77.705 189.210 77.875 189.560 ;
        RECT 67.455 188.980 77.490 189.150 ;
        RECT 67.455 188.420 77.490 188.590 ;
        RECT 67.070 188.010 67.240 188.360 ;
        RECT 77.705 188.010 77.875 188.360 ;
        RECT 67.455 187.780 77.490 187.950 ;
        RECT 76.730 187.390 77.450 187.480 ;
        RECT 67.455 187.220 77.490 187.390 ;
        RECT 67.070 186.810 67.240 187.160 ;
        RECT 76.730 187.140 77.450 187.220 ;
        RECT 77.705 186.810 77.875 187.160 ;
        RECT 67.455 186.580 77.490 186.750 ;
        RECT 78.065 186.250 79.420 191.320 ;
        RECT 85.360 191.390 87.110 191.560 ;
        RECT 85.360 187.900 85.530 191.390 ;
        RECT 86.070 190.880 86.400 191.050 ;
        RECT 85.930 188.625 86.100 190.665 ;
        RECT 86.370 188.625 86.540 190.665 ;
        RECT 86.070 188.240 86.400 188.410 ;
        RECT 86.940 187.900 87.110 191.390 ;
        RECT 85.360 187.730 87.110 187.900 ;
        RECT 87.460 191.390 89.210 191.560 ;
        RECT 87.460 187.900 87.630 191.390 ;
        RECT 88.170 190.880 88.500 191.050 ;
        RECT 88.030 188.625 88.200 190.665 ;
        RECT 88.470 188.625 88.640 190.665 ;
        RECT 88.170 188.240 88.500 188.410 ;
        RECT 89.040 187.900 89.210 191.390 ;
        RECT 87.460 187.730 89.210 187.900 ;
        RECT 85.380 187.690 87.080 187.730 ;
        RECT 87.480 187.690 89.180 187.730 ;
        RECT 85.380 187.370 87.080 187.410 ;
        RECT 87.480 187.370 89.180 187.410 ;
        RECT 54.160 185.170 79.420 186.250 ;
        RECT 54.160 182.910 61.160 185.170 ;
        RECT 61.885 184.600 71.925 184.770 ;
        RECT 61.500 183.540 61.670 184.540 ;
        RECT 72.140 183.540 72.310 184.540 ;
        RECT 61.885 183.310 71.925 183.480 ;
        RECT 61.965 182.910 71.845 183.310 ;
        RECT 72.640 182.910 79.420 185.170 ;
        RECT 85.360 187.200 87.110 187.370 ;
        RECT 85.360 183.710 85.530 187.200 ;
        RECT 86.070 186.690 86.400 186.860 ;
        RECT 85.930 184.435 86.100 186.475 ;
        RECT 86.370 184.435 86.540 186.475 ;
        RECT 86.070 184.050 86.400 184.220 ;
        RECT 86.940 183.710 87.110 187.200 ;
        RECT 85.360 183.540 87.110 183.710 ;
        RECT 87.460 187.200 89.210 187.370 ;
        RECT 87.460 183.710 87.630 187.200 ;
        RECT 88.170 186.690 88.500 186.860 ;
        RECT 88.030 184.435 88.200 186.475 ;
        RECT 88.470 184.435 88.640 186.475 ;
        RECT 88.170 184.050 88.500 184.220 ;
        RECT 89.040 183.710 89.210 187.200 ;
        RECT 87.460 183.540 89.210 183.710 ;
        RECT 54.160 182.300 79.420 182.910 ;
        RECT 54.160 180.040 57.230 182.300 ;
        RECT 57.945 181.730 65.985 181.900 ;
        RECT 57.560 180.670 57.730 181.670 ;
        RECT 66.200 180.670 66.370 181.670 ;
        RECT 57.945 180.440 65.985 180.610 ;
        RECT 66.710 180.040 66.880 182.300 ;
        RECT 72.640 182.290 79.420 182.300 ;
        RECT 67.605 181.730 75.645 181.900 ;
        RECT 67.220 180.670 67.390 181.670 ;
        RECT 75.860 180.670 76.030 181.670 ;
        RECT 67.605 180.440 75.645 180.610 ;
        RECT 76.370 180.040 79.420 182.290 ;
        RECT 85.360 183.010 87.110 183.180 ;
        RECT 85.360 180.610 85.530 183.010 ;
        RECT 86.070 182.500 86.400 182.670 ;
        RECT 85.930 181.290 86.100 182.330 ;
        RECT 86.370 181.290 86.540 182.330 ;
        RECT 86.070 180.950 86.400 181.120 ;
        RECT 86.940 180.610 87.110 183.010 ;
        RECT 85.360 180.440 87.110 180.610 ;
        RECT 87.460 183.010 89.210 183.180 ;
        RECT 87.460 180.610 87.630 183.010 ;
        RECT 88.170 182.500 88.500 182.670 ;
        RECT 88.030 181.290 88.200 182.330 ;
        RECT 88.470 181.290 88.640 182.330 ;
        RECT 88.170 180.950 88.500 181.120 ;
        RECT 89.040 180.610 89.210 183.010 ;
        RECT 87.460 180.440 89.210 180.610 ;
        RECT 85.380 180.410 87.080 180.440 ;
        RECT 87.480 180.410 89.180 180.440 ;
        RECT 85.380 180.080 87.080 180.110 ;
        RECT 87.480 180.080 89.180 180.110 ;
        RECT 54.160 179.870 79.420 180.040 ;
        RECT 85.360 179.910 87.110 180.080 ;
        RECT 12.120 178.830 23.310 179.000 ;
        RECT 12.120 172.140 12.290 178.830 ;
        RECT 12.770 172.620 14.930 178.350 ;
        RECT 20.500 172.620 22.660 178.350 ;
        RECT 23.140 172.140 23.310 178.830 ;
        RECT 12.120 171.970 23.310 172.140 ;
        RECT 12.120 165.280 12.290 171.970 ;
        RECT 12.770 165.760 14.930 171.490 ;
        RECT 20.500 165.760 22.660 171.490 ;
        RECT 23.140 165.280 23.310 171.970 ;
        RECT 27.240 179.340 52.500 179.510 ;
        RECT 27.240 177.080 30.310 179.340 ;
        RECT 31.025 178.770 39.065 178.940 ;
        RECT 30.640 177.710 30.810 178.710 ;
        RECT 39.280 177.710 39.450 178.710 ;
        RECT 31.025 177.480 39.065 177.650 ;
        RECT 39.790 177.080 39.960 179.340 ;
        RECT 40.685 178.770 48.725 178.940 ;
        RECT 40.300 177.710 40.470 178.710 ;
        RECT 48.940 177.710 49.110 178.710 ;
        RECT 40.685 177.480 48.725 177.650 ;
        RECT 49.450 177.090 52.500 179.340 ;
        RECT 45.720 177.080 52.500 177.090 ;
        RECT 27.240 176.470 52.500 177.080 ;
        RECT 27.240 174.210 34.240 176.470 ;
        RECT 35.045 176.070 44.925 176.470 ;
        RECT 34.965 175.900 45.005 176.070 ;
        RECT 34.580 174.840 34.750 175.840 ;
        RECT 45.220 174.840 45.390 175.840 ;
        RECT 34.965 174.610 45.005 174.780 ;
        RECT 45.720 174.210 52.500 176.470 ;
        RECT 27.240 173.130 52.500 174.210 ;
        RECT 27.240 168.060 28.600 173.130 ;
        RECT 29.175 172.630 39.210 172.800 ;
        RECT 28.790 172.220 28.960 172.570 ;
        RECT 39.425 172.220 39.595 172.570 ;
        RECT 29.175 171.990 39.210 172.160 ;
        RECT 29.175 171.430 39.210 171.600 ;
        RECT 28.790 171.020 28.960 171.370 ;
        RECT 39.425 171.020 39.595 171.370 ;
        RECT 29.175 170.790 39.210 170.960 ;
        RECT 29.175 170.230 39.210 170.400 ;
        RECT 28.790 169.820 28.960 170.170 ;
        RECT 39.425 169.820 39.595 170.170 ;
        RECT 29.175 169.590 39.210 169.760 ;
        RECT 29.175 169.030 39.210 169.200 ;
        RECT 28.790 168.620 28.960 168.970 ;
        RECT 39.425 168.620 39.595 168.970 ;
        RECT 29.175 168.390 39.210 168.560 ;
        RECT 39.790 168.060 39.960 173.130 ;
        RECT 40.535 172.630 50.570 172.800 ;
        RECT 40.150 172.220 40.320 172.570 ;
        RECT 49.810 172.160 50.530 172.240 ;
        RECT 50.785 172.220 50.955 172.570 ;
        RECT 40.535 171.990 50.570 172.160 ;
        RECT 49.810 171.900 50.530 171.990 ;
        RECT 40.535 171.430 50.570 171.600 ;
        RECT 40.150 171.020 40.320 171.370 ;
        RECT 50.785 171.020 50.955 171.370 ;
        RECT 40.535 170.790 50.570 170.960 ;
        RECT 40.535 170.230 50.570 170.400 ;
        RECT 40.150 169.820 40.320 170.170 ;
        RECT 49.810 169.760 50.530 169.840 ;
        RECT 50.785 169.820 50.955 170.170 ;
        RECT 40.535 169.590 50.570 169.760 ;
        RECT 49.810 169.500 50.530 169.590 ;
        RECT 40.535 169.030 50.570 169.200 ;
        RECT 40.150 168.620 40.320 168.970 ;
        RECT 50.785 168.620 50.955 168.970 ;
        RECT 40.535 168.390 50.570 168.560 ;
        RECT 51.145 168.060 52.500 173.130 ;
        RECT 27.240 167.890 52.500 168.060 ;
        RECT 54.160 179.340 79.420 179.510 ;
        RECT 54.160 177.080 57.230 179.340 ;
        RECT 57.945 178.770 65.985 178.940 ;
        RECT 57.560 177.710 57.730 178.710 ;
        RECT 66.200 177.710 66.370 178.710 ;
        RECT 57.945 177.480 65.985 177.650 ;
        RECT 66.710 177.080 66.880 179.340 ;
        RECT 67.605 178.770 75.645 178.940 ;
        RECT 67.220 177.710 67.390 178.710 ;
        RECT 75.860 177.710 76.030 178.710 ;
        RECT 67.605 177.480 75.645 177.650 ;
        RECT 76.370 177.090 79.420 179.340 ;
        RECT 85.360 177.510 85.530 179.910 ;
        RECT 86.070 179.400 86.400 179.570 ;
        RECT 85.930 178.190 86.100 179.230 ;
        RECT 86.370 178.190 86.540 179.230 ;
        RECT 86.070 177.850 86.400 178.020 ;
        RECT 86.940 177.510 87.110 179.910 ;
        RECT 85.360 177.340 87.110 177.510 ;
        RECT 87.460 179.910 89.210 180.080 ;
        RECT 87.460 177.510 87.630 179.910 ;
        RECT 88.170 179.400 88.500 179.570 ;
        RECT 88.030 178.190 88.200 179.230 ;
        RECT 88.470 178.190 88.640 179.230 ;
        RECT 88.170 177.850 88.500 178.020 ;
        RECT 89.040 177.510 89.210 179.910 ;
        RECT 87.460 177.340 89.210 177.510 ;
        RECT 72.640 177.080 79.420 177.090 ;
        RECT 54.160 176.470 79.420 177.080 ;
        RECT 54.160 174.210 61.160 176.470 ;
        RECT 61.965 176.070 71.845 176.470 ;
        RECT 61.885 175.900 71.925 176.070 ;
        RECT 61.500 174.840 61.670 175.840 ;
        RECT 72.140 174.840 72.310 175.840 ;
        RECT 61.885 174.610 71.925 174.780 ;
        RECT 72.640 174.210 79.420 176.470 ;
        RECT 54.160 173.130 79.420 174.210 ;
        RECT 85.360 176.810 87.110 176.980 ;
        RECT 85.360 173.320 85.530 176.810 ;
        RECT 86.070 176.300 86.400 176.470 ;
        RECT 85.930 174.045 86.100 176.085 ;
        RECT 86.370 174.045 86.540 176.085 ;
        RECT 86.070 173.660 86.400 173.830 ;
        RECT 86.940 173.320 87.110 176.810 ;
        RECT 85.360 173.150 87.110 173.320 ;
        RECT 87.460 176.810 89.210 176.980 ;
        RECT 87.460 173.320 87.630 176.810 ;
        RECT 88.170 176.300 88.500 176.470 ;
        RECT 88.030 174.045 88.200 176.085 ;
        RECT 88.470 174.045 88.640 176.085 ;
        RECT 88.170 173.660 88.500 173.830 ;
        RECT 89.040 173.320 89.210 176.810 ;
        RECT 87.460 173.150 89.210 173.320 ;
        RECT 54.160 168.060 55.520 173.130 ;
        RECT 56.095 172.630 66.130 172.800 ;
        RECT 55.710 172.220 55.880 172.570 ;
        RECT 66.345 172.220 66.515 172.570 ;
        RECT 56.095 171.990 66.130 172.160 ;
        RECT 56.095 171.430 66.130 171.600 ;
        RECT 55.710 171.020 55.880 171.370 ;
        RECT 66.345 171.020 66.515 171.370 ;
        RECT 56.095 170.790 66.130 170.960 ;
        RECT 56.095 170.230 66.130 170.400 ;
        RECT 55.710 169.820 55.880 170.170 ;
        RECT 66.345 169.820 66.515 170.170 ;
        RECT 56.095 169.590 66.130 169.760 ;
        RECT 56.095 169.030 66.130 169.200 ;
        RECT 55.710 168.620 55.880 168.970 ;
        RECT 66.345 168.620 66.515 168.970 ;
        RECT 56.095 168.390 66.130 168.560 ;
        RECT 66.710 168.060 66.880 173.130 ;
        RECT 67.455 172.630 77.490 172.800 ;
        RECT 67.070 172.220 67.240 172.570 ;
        RECT 76.730 172.160 77.450 172.240 ;
        RECT 77.705 172.220 77.875 172.570 ;
        RECT 67.455 171.990 77.490 172.160 ;
        RECT 76.730 171.900 77.450 171.990 ;
        RECT 67.455 171.430 77.490 171.600 ;
        RECT 67.070 171.020 67.240 171.370 ;
        RECT 77.705 171.020 77.875 171.370 ;
        RECT 67.455 170.790 77.490 170.960 ;
        RECT 67.455 170.230 77.490 170.400 ;
        RECT 67.070 169.820 67.240 170.170 ;
        RECT 76.730 169.760 77.450 169.840 ;
        RECT 77.705 169.820 77.875 170.170 ;
        RECT 67.455 169.590 77.490 169.760 ;
        RECT 76.730 169.500 77.450 169.590 ;
        RECT 67.455 169.030 77.490 169.200 ;
        RECT 67.070 168.620 67.240 168.970 ;
        RECT 77.705 168.620 77.875 168.970 ;
        RECT 67.455 168.390 77.490 168.560 ;
        RECT 78.065 168.060 79.420 173.130 ;
        RECT 85.380 173.110 87.080 173.150 ;
        RECT 87.480 173.110 89.180 173.150 ;
        RECT 85.380 172.790 87.080 172.830 ;
        RECT 87.480 172.790 89.180 172.830 ;
        RECT 85.360 172.620 87.110 172.790 ;
        RECT 85.360 169.130 85.530 172.620 ;
        RECT 86.070 172.110 86.400 172.280 ;
        RECT 85.930 169.855 86.100 171.895 ;
        RECT 86.370 169.855 86.540 171.895 ;
        RECT 86.070 169.470 86.400 169.640 ;
        RECT 86.940 169.130 87.110 172.620 ;
        RECT 85.360 168.960 87.110 169.130 ;
        RECT 87.460 172.620 89.210 172.790 ;
        RECT 87.460 169.130 87.630 172.620 ;
        RECT 88.170 172.110 88.500 172.280 ;
        RECT 88.030 169.855 88.200 171.895 ;
        RECT 88.470 169.855 88.640 171.895 ;
        RECT 88.170 169.470 88.500 169.640 ;
        RECT 89.040 169.130 89.210 172.620 ;
        RECT 87.460 168.960 89.210 169.130 ;
        RECT 54.160 167.890 79.420 168.060 ;
        RECT 85.360 168.430 87.110 168.600 ;
        RECT 12.120 165.110 23.310 165.280 ;
        RECT 12.120 158.420 12.290 165.110 ;
        RECT 12.770 158.900 14.930 164.630 ;
        RECT 20.500 158.900 22.660 164.630 ;
        RECT 23.140 158.420 23.310 165.110 ;
        RECT 27.250 166.220 52.500 166.390 ;
        RECT 27.250 164.370 27.420 166.220 ;
        RECT 28.100 165.650 32.140 165.820 ;
        RECT 27.760 164.590 27.930 165.590 ;
        RECT 32.310 164.590 32.480 165.590 ;
        RECT 28.180 164.530 32.060 164.560 ;
        RECT 28.100 164.370 32.140 164.530 ;
        RECT 32.820 164.370 32.990 166.220 ;
        RECT 33.950 165.650 38.990 165.820 ;
        RECT 33.610 164.590 33.780 165.590 ;
        RECT 39.160 164.590 39.330 165.590 ;
        RECT 33.950 164.370 38.990 164.530 ;
        RECT 39.790 164.370 39.960 166.220 ;
        RECT 40.920 165.650 45.960 165.820 ;
        RECT 40.580 164.590 40.750 165.590 ;
        RECT 46.130 164.590 46.300 165.590 ;
        RECT 40.920 164.370 45.960 164.530 ;
        RECT 46.760 164.370 46.930 166.220 ;
        RECT 47.610 165.650 51.650 165.820 ;
        RECT 47.270 164.590 47.440 165.590 ;
        RECT 51.820 164.590 51.990 165.590 ;
        RECT 47.690 164.530 51.570 164.560 ;
        RECT 47.610 164.370 51.650 164.530 ;
        RECT 52.330 164.370 52.500 166.220 ;
        RECT 54.170 166.220 79.420 166.390 ;
        RECT 54.170 164.370 54.340 166.220 ;
        RECT 55.020 165.650 59.060 165.820 ;
        RECT 54.680 164.590 54.850 165.590 ;
        RECT 59.230 164.590 59.400 165.590 ;
        RECT 55.100 164.530 58.980 164.560 ;
        RECT 55.020 164.370 59.060 164.530 ;
        RECT 59.740 164.370 59.910 166.220 ;
        RECT 60.870 165.650 65.910 165.820 ;
        RECT 60.530 164.590 60.700 165.590 ;
        RECT 66.080 164.590 66.250 165.590 ;
        RECT 60.870 164.370 65.910 164.530 ;
        RECT 66.710 164.370 66.880 166.220 ;
        RECT 67.840 165.650 72.880 165.820 ;
        RECT 67.500 164.590 67.670 165.590 ;
        RECT 73.050 164.590 73.220 165.590 ;
        RECT 67.840 164.370 72.880 164.530 ;
        RECT 73.680 164.370 73.850 166.220 ;
        RECT 74.530 165.650 78.570 165.820 ;
        RECT 74.190 164.590 74.360 165.590 ;
        RECT 78.740 164.590 78.910 165.590 ;
        RECT 74.610 164.530 78.490 164.560 ;
        RECT 74.530 164.370 78.570 164.530 ;
        RECT 79.250 164.370 79.420 166.220 ;
        RECT 85.360 166.030 85.530 168.430 ;
        RECT 86.070 167.920 86.400 168.090 ;
        RECT 85.930 166.710 86.100 167.750 ;
        RECT 86.370 166.710 86.540 167.750 ;
        RECT 86.070 166.370 86.400 166.540 ;
        RECT 86.940 166.030 87.110 168.430 ;
        RECT 85.360 165.860 87.110 166.030 ;
        RECT 87.460 168.430 89.210 168.600 ;
        RECT 87.460 166.030 87.630 168.430 ;
        RECT 88.170 167.920 88.500 168.090 ;
        RECT 88.030 166.710 88.200 167.750 ;
        RECT 88.470 166.710 88.640 167.750 ;
        RECT 88.170 166.370 88.500 166.540 ;
        RECT 89.040 166.030 89.210 168.430 ;
        RECT 87.460 165.860 89.210 166.030 ;
        RECT 85.380 165.830 87.080 165.860 ;
        RECT 87.480 165.830 89.180 165.860 ;
        RECT 27.240 163.790 52.500 164.370 ;
        RECT 27.240 161.530 32.990 163.790 ;
        RECT 33.950 163.220 38.990 163.390 ;
        RECT 33.610 162.160 33.780 163.160 ;
        RECT 39.160 162.160 39.330 163.160 ;
        RECT 33.950 161.930 38.990 162.100 ;
        RECT 39.790 161.530 39.960 163.790 ;
        RECT 40.920 163.220 45.960 163.390 ;
        RECT 40.580 162.160 40.750 163.160 ;
        RECT 46.130 162.160 46.300 163.160 ;
        RECT 40.920 161.930 45.960 162.100 ;
        RECT 46.760 161.530 52.500 163.790 ;
        RECT 27.240 161.360 52.500 161.530 ;
        RECT 54.160 163.790 79.420 164.370 ;
        RECT 54.160 161.530 59.910 163.790 ;
        RECT 60.870 163.220 65.910 163.390 ;
        RECT 60.530 162.160 60.700 163.160 ;
        RECT 66.080 162.160 66.250 163.160 ;
        RECT 60.870 161.930 65.910 162.100 ;
        RECT 66.710 161.530 66.880 163.790 ;
        RECT 67.840 163.220 72.880 163.390 ;
        RECT 67.500 162.160 67.670 163.160 ;
        RECT 73.050 162.160 73.220 163.160 ;
        RECT 67.840 161.930 72.880 162.100 ;
        RECT 73.680 161.530 79.420 163.790 ;
        RECT 54.160 161.360 79.420 161.530 ;
        RECT 54.160 160.830 79.420 161.000 ;
        RECT 44.020 159.660 50.440 159.700 ;
        RECT 12.120 158.250 23.310 158.420 ;
        RECT 12.120 151.560 12.290 158.250 ;
        RECT 12.770 152.040 14.930 157.770 ;
        RECT 20.500 152.040 22.660 157.770 ;
        RECT 23.140 151.560 23.310 158.250 ;
        RECT 43.880 159.490 50.620 159.660 ;
        RECT 43.880 157.230 44.050 159.490 ;
        RECT 44.730 158.920 49.770 159.090 ;
        RECT 44.390 157.860 44.560 158.860 ;
        RECT 49.940 157.860 50.110 158.860 ;
        RECT 44.730 157.630 49.770 157.800 ;
        RECT 50.450 157.230 50.620 159.490 ;
        RECT 54.160 158.570 59.910 160.830 ;
        RECT 60.870 160.260 65.910 160.430 ;
        RECT 60.530 159.200 60.700 160.200 ;
        RECT 66.080 159.200 66.250 160.200 ;
        RECT 60.870 158.970 65.910 159.140 ;
        RECT 66.710 158.570 66.880 160.830 ;
        RECT 67.840 160.260 72.880 160.430 ;
        RECT 67.500 159.200 67.670 160.200 ;
        RECT 73.050 159.200 73.220 160.200 ;
        RECT 67.840 158.970 72.880 159.140 ;
        RECT 73.680 158.570 79.420 160.830 ;
        RECT 54.160 157.990 79.420 158.570 ;
        RECT 43.880 157.060 50.620 157.230 ;
        RECT 44.040 156.785 50.500 157.060 ;
        RECT 12.120 151.390 23.310 151.560 ;
        RECT 12.120 144.700 12.290 151.390 ;
        RECT 12.770 145.180 14.930 150.910 ;
        RECT 20.500 145.180 22.660 150.910 ;
        RECT 23.140 144.700 23.310 151.390 ;
        RECT 38.160 156.615 50.620 156.785 ;
        RECT 38.160 154.255 38.330 156.615 ;
        RECT 38.810 154.735 40.970 156.135 ;
        RECT 47.810 154.735 49.970 156.135 ;
        RECT 50.450 154.255 50.620 156.615 ;
        RECT 54.170 156.140 54.340 157.990 ;
        RECT 55.020 157.830 59.060 157.990 ;
        RECT 55.100 157.800 58.980 157.830 ;
        RECT 54.680 156.770 54.850 157.770 ;
        RECT 59.230 156.770 59.400 157.770 ;
        RECT 55.020 156.540 59.060 156.710 ;
        RECT 59.740 156.140 59.910 157.990 ;
        RECT 60.870 157.830 65.910 157.990 ;
        RECT 60.530 156.770 60.700 157.770 ;
        RECT 66.080 156.770 66.250 157.770 ;
        RECT 60.870 156.540 65.910 156.710 ;
        RECT 66.710 156.140 66.880 157.990 ;
        RECT 67.840 157.830 72.880 157.990 ;
        RECT 67.500 156.770 67.670 157.770 ;
        RECT 73.050 156.770 73.220 157.770 ;
        RECT 67.840 156.540 72.880 156.710 ;
        RECT 73.680 156.140 73.850 157.990 ;
        RECT 74.530 157.830 78.570 157.990 ;
        RECT 74.610 157.800 78.490 157.830 ;
        RECT 74.190 156.770 74.360 157.770 ;
        RECT 78.740 156.770 78.910 157.770 ;
        RECT 74.530 156.540 78.570 156.710 ;
        RECT 79.250 156.140 79.420 157.990 ;
        RECT 54.170 155.970 79.420 156.140 ;
        RECT 38.160 154.075 50.620 154.255 ;
        RECT 38.160 151.715 38.330 154.075 ;
        RECT 38.810 152.195 40.970 153.595 ;
        RECT 47.810 152.195 49.970 153.595 ;
        RECT 50.450 151.715 50.620 154.075 ;
        RECT 38.160 151.535 50.620 151.715 ;
        RECT 38.160 149.175 38.330 151.535 ;
        RECT 38.810 149.655 40.970 151.055 ;
        RECT 47.810 149.655 49.970 151.055 ;
        RECT 50.450 149.175 50.620 151.535 ;
        RECT 38.160 148.995 50.620 149.175 ;
        RECT 38.160 146.635 38.330 148.995 ;
        RECT 38.810 147.115 40.970 148.515 ;
        RECT 47.810 147.115 49.970 148.515 ;
        RECT 50.450 146.635 50.620 148.995 ;
        RECT 38.160 146.465 50.620 146.635 ;
        RECT 54.160 154.300 79.420 154.470 ;
        RECT 54.160 149.230 55.520 154.300 ;
        RECT 56.095 153.800 66.130 153.970 ;
        RECT 55.710 153.390 55.880 153.740 ;
        RECT 66.345 153.390 66.515 153.740 ;
        RECT 56.095 153.160 66.130 153.330 ;
        RECT 56.095 152.600 66.130 152.770 ;
        RECT 55.710 152.190 55.880 152.540 ;
        RECT 66.345 152.190 66.515 152.540 ;
        RECT 56.095 151.960 66.130 152.130 ;
        RECT 56.095 151.400 66.130 151.570 ;
        RECT 55.710 150.990 55.880 151.340 ;
        RECT 66.345 150.990 66.515 151.340 ;
        RECT 56.095 150.760 66.130 150.930 ;
        RECT 56.095 150.200 66.130 150.370 ;
        RECT 55.710 149.790 55.880 150.140 ;
        RECT 66.345 149.790 66.515 150.140 ;
        RECT 56.095 149.560 66.130 149.730 ;
        RECT 66.710 149.230 66.880 154.300 ;
        RECT 67.455 153.800 77.490 153.970 ;
        RECT 67.070 153.390 67.240 153.740 ;
        RECT 77.705 153.390 77.875 153.740 ;
        RECT 67.455 153.160 77.490 153.330 ;
        RECT 76.730 152.770 77.450 152.860 ;
        RECT 67.455 152.600 77.490 152.770 ;
        RECT 67.070 152.190 67.240 152.540 ;
        RECT 76.730 152.520 77.450 152.600 ;
        RECT 77.705 152.190 77.875 152.540 ;
        RECT 67.455 151.960 77.490 152.130 ;
        RECT 67.455 151.400 77.490 151.570 ;
        RECT 67.070 150.990 67.240 151.340 ;
        RECT 77.705 150.990 77.875 151.340 ;
        RECT 67.455 150.760 77.490 150.930 ;
        RECT 76.730 150.370 77.450 150.460 ;
        RECT 67.455 150.200 77.490 150.370 ;
        RECT 67.070 149.790 67.240 150.140 ;
        RECT 76.730 150.120 77.450 150.200 ;
        RECT 77.705 149.790 77.875 150.140 ;
        RECT 67.455 149.560 77.490 149.730 ;
        RECT 78.065 149.230 79.420 154.300 ;
        RECT 54.160 148.150 79.420 149.230 ;
        RECT 54.160 145.890 61.160 148.150 ;
        RECT 61.885 147.580 71.925 147.750 ;
        RECT 61.500 146.520 61.670 147.520 ;
        RECT 72.140 146.520 72.310 147.520 ;
        RECT 61.885 146.290 71.925 146.460 ;
        RECT 61.965 145.890 71.845 146.290 ;
        RECT 72.640 145.890 79.420 148.150 ;
        RECT 54.160 145.280 79.420 145.890 ;
        RECT 39.425 145.030 49.465 145.200 ;
        RECT 12.120 144.530 23.310 144.700 ;
        RECT 39.035 143.970 39.205 144.970 ;
        RECT 49.685 143.970 49.855 144.970 ;
        RECT 39.425 143.740 49.465 143.910 ;
        RECT 38.690 143.150 50.340 143.340 ;
        RECT 54.160 143.020 57.230 145.280 ;
        RECT 57.945 144.710 65.985 144.880 ;
        RECT 57.560 143.650 57.730 144.650 ;
        RECT 66.200 143.650 66.370 144.650 ;
        RECT 57.945 143.420 65.985 143.590 ;
        RECT 66.710 143.020 66.880 145.280 ;
        RECT 72.640 145.270 79.420 145.280 ;
        RECT 67.605 144.710 75.645 144.880 ;
        RECT 67.220 143.650 67.390 144.650 ;
        RECT 75.860 143.650 76.030 144.650 ;
        RECT 67.605 143.420 75.645 143.590 ;
        RECT 76.370 143.020 79.420 145.270 ;
        RECT 54.160 142.850 79.420 143.020 ;
      LAYER met1 ;
        RECT 27.070 216.330 104.140 217.740 ;
        RECT 11.940 213.030 23.490 215.190 ;
        RECT 27.070 214.100 30.310 216.330 ;
        RECT 31.105 215.990 38.985 216.330 ;
        RECT 40.765 215.990 48.645 216.330 ;
        RECT 31.045 215.760 39.045 215.990 ;
        RECT 40.705 215.760 48.705 215.990 ;
        RECT 30.610 215.370 30.840 215.710 ;
        RECT 39.250 215.650 39.480 215.710 ;
        RECT 40.270 215.650 40.500 215.710 ;
        RECT 39.250 215.370 40.500 215.650 ;
        RECT 48.910 215.370 49.140 215.710 ;
        RECT 30.610 215.110 49.140 215.370 ;
        RECT 30.610 214.720 30.840 215.110 ;
        RECT 39.250 214.810 40.500 215.110 ;
        RECT 39.250 214.720 39.480 214.810 ;
        RECT 40.270 214.750 40.500 214.810 ;
        RECT 48.910 214.750 49.140 215.110 ;
        RECT 30.610 214.460 39.480 214.720 ;
        RECT 40.710 214.700 48.690 214.720 ;
        RECT 40.705 214.470 48.705 214.700 ;
        RECT 40.710 214.460 48.690 214.470 ;
        RECT 49.440 214.100 57.240 216.330 ;
        RECT 58.025 215.990 65.905 216.330 ;
        RECT 67.685 215.990 75.565 216.330 ;
        RECT 76.360 216.310 104.140 216.330 ;
        RECT 57.965 215.760 65.965 215.990 ;
        RECT 67.625 215.760 75.625 215.990 ;
        RECT 57.530 215.370 57.760 215.710 ;
        RECT 66.170 215.650 66.400 215.710 ;
        RECT 67.190 215.650 67.420 215.710 ;
        RECT 66.170 215.370 67.420 215.650 ;
        RECT 75.830 215.370 76.060 215.710 ;
        RECT 57.530 215.110 76.060 215.370 ;
        RECT 57.530 214.720 57.760 215.110 ;
        RECT 66.170 214.810 67.420 215.110 ;
        RECT 66.170 214.720 66.400 214.810 ;
        RECT 67.190 214.750 67.420 214.810 ;
        RECT 75.830 214.750 76.060 215.110 ;
        RECT 57.530 214.460 66.400 214.720 ;
        RECT 67.630 214.700 75.610 214.720 ;
        RECT 67.625 214.470 75.625 214.700 ;
        RECT 67.630 214.460 75.610 214.470 ;
        RECT 76.360 214.100 79.600 216.310 ;
        RECT 27.070 213.740 79.600 214.100 ;
        RECT 85.380 215.520 85.680 216.310 ;
        RECT 86.080 215.820 86.380 216.120 ;
        RECT 85.900 215.520 86.130 215.615 ;
        RECT 85.380 213.620 86.130 215.520 ;
        RECT 85.900 213.615 86.130 213.620 ;
        RECT 86.340 215.520 86.570 215.615 ;
        RECT 87.480 215.520 87.780 216.310 ;
        RECT 88.180 215.820 88.480 216.120 ;
        RECT 88.000 215.520 88.230 215.615 ;
        RECT 86.340 213.620 86.980 215.520 ;
        RECT 87.480 213.620 88.230 215.520 ;
        RECT 86.340 213.615 86.570 213.620 ;
        RECT 12.770 200.060 14.930 213.030 ;
        RECT 34.985 212.890 44.985 213.120 ;
        RECT 34.550 212.780 34.780 212.840 ;
        RECT 45.190 212.780 45.420 212.840 ;
        RECT 12.770 186.340 14.930 198.930 ;
        RECT 20.500 193.200 22.660 212.650 ;
        RECT 34.480 211.940 34.840 212.780 ;
        RECT 45.120 211.940 45.480 212.780 ;
        RECT 34.550 211.880 34.780 211.940 ;
        RECT 45.190 211.880 45.420 211.940 ;
        RECT 34.995 211.830 44.975 211.860 ;
        RECT 34.985 211.600 44.985 211.830 ;
        RECT 24.450 210.760 25.180 211.590 ;
        RECT 51.000 211.570 51.730 213.240 ;
        RECT 61.905 212.890 71.905 213.120 ;
        RECT 61.470 212.780 61.700 212.840 ;
        RECT 72.110 212.780 72.340 212.840 ;
        RECT 61.400 211.940 61.760 212.780 ;
        RECT 72.040 211.940 72.400 212.780 ;
        RECT 79.210 212.720 80.310 212.920 ;
        RECT 84.300 212.720 85.420 213.000 ;
        RECT 86.080 212.720 86.380 213.420 ;
        RECT 79.210 212.320 86.380 212.720 ;
        RECT 79.210 212.110 80.310 212.320 ;
        RECT 84.300 212.030 85.420 212.320 ;
        RECT 61.470 211.880 61.700 211.940 ;
        RECT 72.110 211.880 72.340 211.940 ;
        RECT 61.915 211.830 71.895 211.860 ;
        RECT 61.905 211.600 71.905 211.830 ;
        RECT 86.080 211.620 86.380 212.320 ;
        RECT 86.780 212.720 86.980 213.620 ;
        RECT 88.000 213.615 88.230 213.620 ;
        RECT 88.440 215.520 88.670 215.615 ;
        RECT 89.550 215.560 89.880 216.310 ;
        RECT 90.280 215.820 92.190 216.100 ;
        RECT 93.440 215.830 93.770 216.100 ;
        RECT 93.460 215.820 93.750 215.830 ;
        RECT 90.110 215.560 90.340 215.615 ;
        RECT 88.440 213.620 89.080 215.520 ;
        RECT 89.550 213.670 90.340 215.560 ;
        RECT 88.440 213.615 88.670 213.620 ;
        RECT 88.180 212.720 88.480 213.420 ;
        RECT 86.780 212.320 88.480 212.720 ;
        RECT 51.000 211.210 54.410 211.570 ;
        RECT 85.900 211.420 86.130 211.470 ;
        RECT 53.990 210.760 54.410 211.210 ;
        RECT 24.450 210.500 51.370 210.760 ;
        RECT 53.990 210.500 78.290 210.760 ;
        RECT 24.450 209.560 25.180 210.500 ;
        RECT 38.480 209.850 39.200 209.890 ;
        RECT 40.560 209.850 41.260 209.860 ;
        RECT 29.195 209.620 39.200 209.850 ;
        RECT 40.555 209.620 50.550 209.850 ;
        RECT 38.480 209.570 39.200 209.620 ;
        RECT 40.560 209.590 41.650 209.620 ;
        RECT 28.740 209.510 29.020 209.570 ;
        RECT 28.390 209.320 29.020 209.510 ;
        RECT 28.390 207.110 28.580 209.320 ;
        RECT 28.740 209.260 29.020 209.320 ;
        RECT 39.380 209.260 39.650 209.570 ;
        RECT 40.100 209.260 40.380 209.570 ;
        RECT 50.740 209.510 51.010 209.570 ;
        RECT 51.180 209.510 51.370 210.500 ;
        RECT 65.400 209.850 66.120 209.890 ;
        RECT 67.480 209.850 68.180 209.860 ;
        RECT 56.115 209.620 66.120 209.850 ;
        RECT 67.475 209.620 77.470 209.850 ;
        RECT 65.400 209.570 66.120 209.620 ;
        RECT 67.480 209.590 68.570 209.620 ;
        RECT 55.660 209.510 55.940 209.570 ;
        RECT 50.740 209.320 51.370 209.510 ;
        RECT 50.740 209.260 51.010 209.320 ;
        RECT 29.220 209.210 29.940 209.250 ;
        RECT 40.550 209.210 41.650 209.220 ;
        RECT 49.810 209.210 50.530 209.260 ;
        RECT 29.195 208.980 39.190 209.210 ;
        RECT 40.550 208.980 50.550 209.210 ;
        RECT 29.220 208.930 29.940 208.980 ;
        RECT 40.550 208.960 41.650 208.980 ;
        RECT 49.810 208.920 50.530 208.980 ;
        RECT 38.480 208.650 39.200 208.690 ;
        RECT 40.560 208.650 41.280 208.700 ;
        RECT 29.195 208.420 39.200 208.650 ;
        RECT 40.555 208.420 50.550 208.650 ;
        RECT 38.480 208.370 39.200 208.420 ;
        RECT 28.720 208.060 29.040 208.370 ;
        RECT 39.340 208.040 39.680 208.390 ;
        RECT 40.070 208.040 40.410 208.390 ;
        RECT 40.560 208.370 41.280 208.420 ;
        RECT 50.710 208.040 51.040 208.400 ;
        RECT 30.420 208.010 31.140 208.040 ;
        RECT 48.610 208.010 49.330 208.020 ;
        RECT 29.195 207.780 39.190 208.010 ;
        RECT 40.555 207.780 50.550 208.010 ;
        RECT 30.420 207.730 31.140 207.780 ;
        RECT 48.610 207.760 49.330 207.780 ;
        RECT 38.480 207.450 39.200 207.490 ;
        RECT 40.560 207.450 41.280 207.500 ;
        RECT 29.195 207.220 39.200 207.450 ;
        RECT 40.555 207.220 50.550 207.450 ;
        RECT 38.480 207.170 39.200 207.220 ;
        RECT 40.560 207.190 41.610 207.220 ;
        RECT 28.740 207.110 29.020 207.170 ;
        RECT 28.390 206.920 29.020 207.110 ;
        RECT 28.390 204.810 28.580 206.920 ;
        RECT 28.740 206.860 29.020 206.920 ;
        RECT 39.380 206.860 39.650 207.170 ;
        RECT 40.100 206.860 40.380 207.170 ;
        RECT 50.740 207.110 51.010 207.170 ;
        RECT 51.180 207.110 51.370 209.320 ;
        RECT 50.740 206.920 51.370 207.110 ;
        RECT 55.310 209.320 55.940 209.510 ;
        RECT 55.310 207.110 55.500 209.320 ;
        RECT 55.660 209.260 55.940 209.320 ;
        RECT 66.300 209.260 66.570 209.570 ;
        RECT 67.020 209.260 67.300 209.570 ;
        RECT 77.660 209.510 77.930 209.570 ;
        RECT 78.100 209.510 78.290 210.500 ;
        RECT 85.380 210.520 86.130 211.420 ;
        RECT 85.380 209.820 85.680 210.520 ;
        RECT 85.900 210.470 86.130 210.520 ;
        RECT 86.340 211.420 86.570 211.470 ;
        RECT 86.780 211.420 86.980 212.320 ;
        RECT 88.180 211.620 88.480 212.320 ;
        RECT 88.880 212.720 89.080 213.620 ;
        RECT 90.110 213.615 90.340 213.670 ;
        RECT 90.550 215.560 90.780 215.615 ;
        RECT 91.690 215.560 91.920 215.615 ;
        RECT 90.550 213.680 91.190 215.560 ;
        RECT 90.550 213.615 90.780 213.680 ;
        RECT 90.300 213.400 90.590 213.410 ;
        RECT 88.880 212.320 89.280 212.720 ;
        RECT 88.000 211.420 88.230 211.470 ;
        RECT 86.340 210.520 86.980 211.420 ;
        RECT 87.480 210.520 88.230 211.420 ;
        RECT 86.340 210.470 86.570 210.520 ;
        RECT 86.080 210.020 86.380 210.320 ;
        RECT 87.480 209.820 87.780 210.520 ;
        RECT 88.000 210.470 88.230 210.520 ;
        RECT 88.440 211.420 88.670 211.470 ;
        RECT 88.880 211.420 89.080 212.320 ;
        RECT 90.280 211.640 90.610 213.400 ;
        RECT 90.930 212.690 91.190 213.680 ;
        RECT 91.370 213.680 91.920 215.560 ;
        RECT 90.900 212.340 91.230 212.690 ;
        RECT 90.300 211.630 90.590 211.640 ;
        RECT 88.440 210.520 89.080 211.420 ;
        RECT 90.110 211.410 90.340 211.470 ;
        RECT 89.520 210.530 90.340 211.410 ;
        RECT 88.440 210.470 88.670 210.520 ;
        RECT 88.180 210.020 88.480 210.320 ;
        RECT 89.520 209.820 89.810 210.530 ;
        RECT 90.110 210.470 90.340 210.530 ;
        RECT 90.550 211.410 90.780 211.470 ;
        RECT 90.930 211.410 91.190 212.340 ;
        RECT 90.550 210.530 91.190 211.410 ;
        RECT 91.370 211.410 91.550 213.680 ;
        RECT 91.690 213.615 91.920 213.680 ;
        RECT 92.130 215.560 92.360 215.615 ;
        RECT 93.270 215.560 93.500 215.615 ;
        RECT 92.130 213.670 93.500 215.560 ;
        RECT 92.130 213.615 92.360 213.670 ;
        RECT 91.860 213.130 92.190 213.410 ;
        RECT 91.860 211.630 92.190 212.680 ;
        RECT 91.690 211.410 91.920 211.470 ;
        RECT 91.370 210.530 91.920 211.410 ;
        RECT 90.550 210.470 90.780 210.530 ;
        RECT 91.690 210.470 91.920 210.530 ;
        RECT 92.130 211.410 92.360 211.470 ;
        RECT 92.500 211.410 93.130 213.670 ;
        RECT 93.270 213.615 93.500 213.670 ;
        RECT 93.710 215.560 93.940 215.615 ;
        RECT 93.710 213.670 94.360 215.560 ;
        RECT 93.710 213.615 93.940 213.670 ;
        RECT 93.440 212.360 93.770 213.410 ;
        RECT 93.440 211.650 93.770 211.910 ;
        RECT 93.460 211.630 93.750 211.650 ;
        RECT 93.270 211.410 93.500 211.470 ;
        RECT 92.130 210.530 93.500 211.410 ;
        RECT 92.130 210.470 92.360 210.530 ;
        RECT 93.270 210.470 93.500 210.530 ;
        RECT 93.710 211.410 93.940 211.470 ;
        RECT 94.080 211.410 94.360 213.670 ;
        RECT 100.130 215.520 100.430 216.310 ;
        RECT 100.830 215.820 101.130 216.120 ;
        RECT 100.650 215.520 100.880 215.615 ;
        RECT 100.130 213.620 100.880 215.520 ;
        RECT 100.650 213.615 100.880 213.620 ;
        RECT 101.090 215.520 101.320 215.615 ;
        RECT 102.230 215.520 102.530 216.310 ;
        RECT 102.930 215.820 103.230 216.120 ;
        RECT 102.750 215.520 102.980 215.615 ;
        RECT 101.090 213.620 101.730 215.520 ;
        RECT 102.230 213.620 102.980 215.520 ;
        RECT 101.090 213.615 101.320 213.620 ;
        RECT 100.830 212.720 101.130 213.420 ;
        RECT 100.130 212.320 101.130 212.720 ;
        RECT 100.830 211.620 101.130 212.320 ;
        RECT 101.530 212.720 101.730 213.620 ;
        RECT 102.750 213.615 102.980 213.620 ;
        RECT 103.190 215.520 103.420 215.615 ;
        RECT 103.190 213.620 103.830 215.520 ;
        RECT 103.190 213.615 103.420 213.620 ;
        RECT 102.930 212.720 103.230 213.420 ;
        RECT 101.530 212.320 103.230 212.720 ;
        RECT 100.650 211.420 100.880 211.470 ;
        RECT 93.710 210.530 94.360 211.410 ;
        RECT 93.710 210.470 93.940 210.530 ;
        RECT 100.130 210.520 100.880 211.420 ;
        RECT 90.300 210.300 90.590 210.310 ;
        RECT 91.880 210.300 92.170 210.310 ;
        RECT 93.460 210.300 93.750 210.310 ;
        RECT 90.180 209.970 90.710 210.300 ;
        RECT 91.860 210.030 92.190 210.300 ;
        RECT 93.330 209.970 93.860 210.300 ;
        RECT 100.130 209.820 100.430 210.520 ;
        RECT 100.650 210.470 100.880 210.520 ;
        RECT 101.090 211.420 101.320 211.470 ;
        RECT 101.530 211.420 101.730 212.320 ;
        RECT 102.930 211.620 103.230 212.320 ;
        RECT 103.630 212.720 103.830 213.620 ;
        RECT 104.630 212.720 105.100 213.490 ;
        RECT 103.630 212.320 105.100 212.720 ;
        RECT 102.750 211.420 102.980 211.470 ;
        RECT 101.090 210.520 101.730 211.420 ;
        RECT 102.230 210.520 102.980 211.420 ;
        RECT 101.090 210.470 101.320 210.520 ;
        RECT 100.830 210.020 101.130 210.320 ;
        RECT 102.230 209.820 102.530 210.520 ;
        RECT 102.750 210.470 102.980 210.520 ;
        RECT 103.190 211.420 103.420 211.470 ;
        RECT 103.630 211.420 103.830 212.320 ;
        RECT 103.190 210.520 103.830 211.420 ;
        RECT 103.190 210.470 103.420 210.520 ;
        RECT 102.930 210.020 103.230 210.320 ;
        RECT 77.660 209.320 78.290 209.510 ;
        RECT 77.660 209.260 77.930 209.320 ;
        RECT 56.140 209.210 56.860 209.250 ;
        RECT 67.470 209.210 68.570 209.220 ;
        RECT 76.730 209.210 77.450 209.260 ;
        RECT 56.115 208.980 66.110 209.210 ;
        RECT 67.470 208.980 77.470 209.210 ;
        RECT 56.140 208.930 56.860 208.980 ;
        RECT 67.470 208.960 68.570 208.980 ;
        RECT 76.730 208.920 77.450 208.980 ;
        RECT 65.400 208.650 66.120 208.690 ;
        RECT 67.480 208.650 68.200 208.700 ;
        RECT 56.115 208.420 66.120 208.650 ;
        RECT 67.475 208.420 77.470 208.650 ;
        RECT 65.400 208.370 66.120 208.420 ;
        RECT 55.640 208.060 55.960 208.370 ;
        RECT 66.260 208.040 66.600 208.390 ;
        RECT 66.990 208.040 67.330 208.390 ;
        RECT 67.480 208.370 68.200 208.420 ;
        RECT 77.630 208.040 77.960 208.400 ;
        RECT 57.340 208.010 58.060 208.040 ;
        RECT 75.530 208.010 76.250 208.020 ;
        RECT 56.115 207.780 66.110 208.010 ;
        RECT 67.475 207.780 77.470 208.010 ;
        RECT 57.340 207.730 58.060 207.780 ;
        RECT 75.530 207.760 76.250 207.780 ;
        RECT 65.400 207.450 66.120 207.490 ;
        RECT 67.480 207.450 68.200 207.500 ;
        RECT 56.115 207.220 66.120 207.450 ;
        RECT 67.475 207.220 77.470 207.450 ;
        RECT 65.400 207.170 66.120 207.220 ;
        RECT 67.480 207.190 68.530 207.220 ;
        RECT 55.660 207.110 55.940 207.170 ;
        RECT 55.310 206.920 55.940 207.110 ;
        RECT 50.740 206.860 51.010 206.920 ;
        RECT 29.220 206.810 29.940 206.850 ;
        RECT 40.550 206.810 41.610 206.820 ;
        RECT 49.810 206.810 50.530 206.860 ;
        RECT 29.195 206.580 39.190 206.810 ;
        RECT 40.550 206.580 50.550 206.810 ;
        RECT 29.220 206.530 29.940 206.580 ;
        RECT 40.550 206.560 41.610 206.580 ;
        RECT 49.810 206.520 50.530 206.580 ;
        RECT 38.480 206.250 39.200 206.290 ;
        RECT 40.560 206.250 41.280 206.300 ;
        RECT 29.195 206.020 39.200 206.250 ;
        RECT 40.555 206.020 50.550 206.250 ;
        RECT 38.480 205.970 39.200 206.020 ;
        RECT 28.720 205.660 29.040 205.970 ;
        RECT 39.340 205.640 39.680 205.990 ;
        RECT 40.070 205.640 40.410 205.990 ;
        RECT 40.560 205.970 41.280 206.020 ;
        RECT 50.710 205.640 51.040 206.000 ;
        RECT 30.420 205.610 31.140 205.640 ;
        RECT 48.610 205.610 49.330 205.620 ;
        RECT 29.195 205.380 39.190 205.610 ;
        RECT 40.555 205.380 50.550 205.610 ;
        RECT 30.420 205.330 31.140 205.380 ;
        RECT 48.610 205.360 49.330 205.380 ;
        RECT 52.970 204.810 53.610 205.830 ;
        RECT 55.310 204.810 55.500 206.920 ;
        RECT 55.660 206.860 55.940 206.920 ;
        RECT 66.300 206.860 66.570 207.170 ;
        RECT 67.020 206.860 67.300 207.170 ;
        RECT 77.660 207.110 77.930 207.170 ;
        RECT 78.100 207.110 78.290 209.320 ;
        RECT 85.180 209.020 104.140 209.820 ;
        RECT 85.380 208.320 85.680 209.020 ;
        RECT 86.080 208.520 86.380 208.820 ;
        RECT 85.900 208.320 86.130 208.370 ;
        RECT 85.380 207.420 86.130 208.320 ;
        RECT 85.900 207.370 86.130 207.420 ;
        RECT 86.340 208.320 86.570 208.370 ;
        RECT 87.480 208.320 87.780 209.020 ;
        RECT 88.180 208.520 88.480 208.820 ;
        RECT 88.000 208.320 88.230 208.370 ;
        RECT 86.340 207.420 86.980 208.320 ;
        RECT 87.480 207.420 88.230 208.320 ;
        RECT 86.340 207.370 86.570 207.420 ;
        RECT 77.660 206.920 78.290 207.110 ;
        RECT 77.660 206.860 77.930 206.920 ;
        RECT 56.140 206.810 56.860 206.850 ;
        RECT 67.470 206.810 68.530 206.820 ;
        RECT 76.730 206.810 77.450 206.860 ;
        RECT 56.115 206.580 66.110 206.810 ;
        RECT 67.470 206.580 77.470 206.810 ;
        RECT 56.140 206.530 56.860 206.580 ;
        RECT 67.470 206.560 68.530 206.580 ;
        RECT 76.730 206.520 77.450 206.580 ;
        RECT 86.080 206.520 86.380 207.220 ;
        RECT 65.400 206.250 66.120 206.290 ;
        RECT 67.480 206.250 68.200 206.300 ;
        RECT 56.115 206.020 66.120 206.250 ;
        RECT 67.475 206.020 77.470 206.250 ;
        RECT 83.140 206.120 86.380 206.520 ;
        RECT 65.400 205.970 66.120 206.020 ;
        RECT 55.640 205.660 55.960 205.970 ;
        RECT 66.260 205.640 66.600 205.990 ;
        RECT 66.990 205.640 67.330 205.990 ;
        RECT 67.480 205.970 68.200 206.020 ;
        RECT 77.630 205.640 77.960 206.000 ;
        RECT 83.140 205.650 84.680 206.120 ;
        RECT 57.340 205.610 58.060 205.640 ;
        RECT 75.530 205.610 76.250 205.620 ;
        RECT 56.115 205.380 66.110 205.610 ;
        RECT 67.475 205.380 77.470 205.610 ;
        RECT 86.080 205.420 86.380 206.120 ;
        RECT 86.780 206.520 86.980 207.420 ;
        RECT 88.000 207.370 88.230 207.420 ;
        RECT 88.440 208.320 88.670 208.370 ;
        RECT 88.440 207.420 89.080 208.320 ;
        RECT 89.520 208.310 89.810 209.020 ;
        RECT 90.180 208.540 90.710 208.870 ;
        RECT 91.860 208.540 92.190 208.810 ;
        RECT 93.330 208.540 93.860 208.870 ;
        RECT 90.300 208.530 90.590 208.540 ;
        RECT 91.880 208.530 92.170 208.540 ;
        RECT 93.460 208.530 93.750 208.540 ;
        RECT 90.110 208.310 90.340 208.370 ;
        RECT 89.520 207.430 90.340 208.310 ;
        RECT 88.440 207.370 88.670 207.420 ;
        RECT 88.180 206.520 88.480 207.220 ;
        RECT 86.780 206.120 88.480 206.520 ;
        RECT 57.340 205.330 58.060 205.380 ;
        RECT 75.530 205.360 76.250 205.380 ;
        RECT 85.900 205.220 86.130 205.225 ;
        RECT 24.620 204.550 51.040 204.810 ;
        RECT 52.970 204.550 77.960 204.810 ;
        RECT 24.620 197.310 25.240 204.550 ;
        RECT 30.410 204.150 50.530 204.410 ;
        RECT 29.210 203.750 49.330 204.010 ;
        RECT 52.970 203.450 53.610 204.550 ;
        RECT 57.330 204.150 77.450 204.410 ;
        RECT 56.130 203.750 76.250 204.010 ;
        RECT 85.380 203.320 86.130 205.220 ;
        RECT 27.730 202.870 32.110 202.890 ;
        RECT 33.980 202.870 38.960 202.890 ;
        RECT 40.950 202.870 45.930 202.890 ;
        RECT 27.730 202.630 32.510 202.870 ;
        RECT 33.970 202.640 38.970 202.870 ;
        RECT 40.940 202.640 45.940 202.870 ;
        RECT 33.980 202.630 38.960 202.640 ;
        RECT 40.950 202.630 45.930 202.640 ;
        RECT 47.270 202.630 52.020 202.890 ;
        RECT 27.730 202.240 27.960 202.630 ;
        RECT 32.280 202.530 32.510 202.630 ;
        RECT 47.270 202.610 47.630 202.630 ;
        RECT 47.270 202.590 47.470 202.610 ;
        RECT 33.580 202.530 33.810 202.590 ;
        RECT 39.130 202.530 39.360 202.590 ;
        RECT 40.550 202.530 40.780 202.590 ;
        RECT 46.100 202.530 46.330 202.590 ;
        RECT 47.240 202.530 47.470 202.590 ;
        RECT 32.280 202.240 33.810 202.530 ;
        RECT 39.060 202.240 39.420 202.530 ;
        RECT 27.730 201.980 39.420 202.240 ;
        RECT 27.730 201.630 27.960 201.980 ;
        RECT 32.280 201.690 33.810 201.980 ;
        RECT 39.060 201.690 39.420 201.980 ;
        RECT 40.490 202.240 40.850 202.530 ;
        RECT 46.100 202.240 47.470 202.530 ;
        RECT 51.790 202.240 52.020 202.630 ;
        RECT 40.490 201.980 52.020 202.240 ;
        RECT 40.490 201.690 40.850 201.980 ;
        RECT 46.100 201.690 47.470 201.980 ;
        RECT 32.280 201.630 32.510 201.690 ;
        RECT 33.580 201.630 33.810 201.690 ;
        RECT 39.130 201.630 39.360 201.690 ;
        RECT 40.550 201.630 40.780 201.690 ;
        RECT 46.100 201.630 46.330 201.690 ;
        RECT 47.240 201.630 47.470 201.690 ;
        RECT 51.790 201.630 52.020 201.980 ;
        RECT 54.650 202.870 59.030 202.890 ;
        RECT 60.900 202.870 65.880 202.890 ;
        RECT 67.870 202.870 72.850 202.890 ;
        RECT 54.650 202.630 59.430 202.870 ;
        RECT 60.890 202.640 65.890 202.870 ;
        RECT 67.860 202.640 72.860 202.870 ;
        RECT 60.900 202.630 65.880 202.640 ;
        RECT 67.870 202.630 72.850 202.640 ;
        RECT 74.190 202.630 78.940 202.890 ;
        RECT 54.650 202.240 54.880 202.630 ;
        RECT 59.200 202.530 59.430 202.630 ;
        RECT 74.190 202.610 74.550 202.630 ;
        RECT 74.190 202.590 74.390 202.610 ;
        RECT 60.500 202.530 60.730 202.590 ;
        RECT 66.050 202.530 66.280 202.590 ;
        RECT 67.470 202.530 67.700 202.590 ;
        RECT 73.020 202.530 73.250 202.590 ;
        RECT 74.160 202.530 74.390 202.590 ;
        RECT 59.200 202.240 60.730 202.530 ;
        RECT 65.980 202.240 66.340 202.530 ;
        RECT 54.650 201.980 66.340 202.240 ;
        RECT 54.650 201.630 54.880 201.980 ;
        RECT 59.200 201.690 60.730 201.980 ;
        RECT 65.980 201.690 66.340 201.980 ;
        RECT 67.410 202.240 67.770 202.530 ;
        RECT 73.020 202.240 74.390 202.530 ;
        RECT 78.710 202.240 78.940 202.630 ;
        RECT 85.380 202.530 85.680 203.320 ;
        RECT 85.900 203.225 86.130 203.320 ;
        RECT 86.340 205.220 86.570 205.225 ;
        RECT 86.780 205.220 86.980 206.120 ;
        RECT 88.180 205.420 88.480 206.120 ;
        RECT 88.880 206.520 89.080 207.420 ;
        RECT 90.110 207.370 90.340 207.430 ;
        RECT 90.550 208.310 90.780 208.370 ;
        RECT 91.690 208.310 91.920 208.370 ;
        RECT 90.550 207.430 91.190 208.310 ;
        RECT 90.550 207.370 90.780 207.430 ;
        RECT 90.300 207.200 90.590 207.210 ;
        RECT 88.880 206.120 89.280 206.520 ;
        RECT 88.000 205.220 88.230 205.225 ;
        RECT 86.340 203.320 86.980 205.220 ;
        RECT 87.480 203.320 88.230 205.220 ;
        RECT 86.340 203.225 86.570 203.320 ;
        RECT 86.080 202.720 86.380 203.020 ;
        RECT 87.480 202.530 87.780 203.320 ;
        RECT 88.000 203.225 88.230 203.320 ;
        RECT 88.440 205.220 88.670 205.225 ;
        RECT 88.880 205.220 89.080 206.120 ;
        RECT 90.280 205.440 90.610 207.200 ;
        RECT 90.930 206.500 91.190 207.430 ;
        RECT 91.370 207.430 91.920 208.310 ;
        RECT 90.900 206.150 91.230 206.500 ;
        RECT 90.300 205.430 90.590 205.440 ;
        RECT 88.440 203.320 89.080 205.220 ;
        RECT 90.110 205.170 90.340 205.225 ;
        RECT 88.440 203.225 88.670 203.320 ;
        RECT 89.550 203.280 90.340 205.170 ;
        RECT 88.180 202.720 88.480 203.020 ;
        RECT 89.550 202.530 89.880 203.280 ;
        RECT 90.110 203.225 90.340 203.280 ;
        RECT 90.550 205.160 90.780 205.225 ;
        RECT 90.930 205.160 91.190 206.150 ;
        RECT 90.550 203.280 91.190 205.160 ;
        RECT 91.370 205.160 91.550 207.430 ;
        RECT 91.690 207.370 91.920 207.430 ;
        RECT 92.130 208.310 92.360 208.370 ;
        RECT 93.270 208.310 93.500 208.370 ;
        RECT 92.130 207.430 93.500 208.310 ;
        RECT 92.130 207.370 92.360 207.430 ;
        RECT 91.860 206.160 92.190 207.210 ;
        RECT 91.860 205.430 92.190 205.710 ;
        RECT 91.690 205.160 91.920 205.225 ;
        RECT 91.370 203.280 91.920 205.160 ;
        RECT 90.550 203.225 90.780 203.280 ;
        RECT 91.690 203.225 91.920 203.280 ;
        RECT 92.130 205.170 92.360 205.225 ;
        RECT 92.500 205.170 93.130 207.430 ;
        RECT 93.270 207.370 93.500 207.430 ;
        RECT 93.710 208.310 93.940 208.370 ;
        RECT 94.790 208.310 95.080 209.020 ;
        RECT 95.450 208.540 95.980 208.870 ;
        RECT 97.130 208.540 97.460 208.810 ;
        RECT 98.600 208.540 99.130 208.870 ;
        RECT 95.570 208.530 95.860 208.540 ;
        RECT 97.150 208.530 97.440 208.540 ;
        RECT 98.730 208.530 99.020 208.540 ;
        RECT 95.380 208.310 95.610 208.370 ;
        RECT 93.710 207.430 94.360 208.310 ;
        RECT 94.790 207.430 95.610 208.310 ;
        RECT 93.710 207.370 93.940 207.430 ;
        RECT 93.460 207.190 93.750 207.210 ;
        RECT 93.440 206.930 93.770 207.190 ;
        RECT 93.440 205.430 93.770 206.480 ;
        RECT 93.270 205.170 93.500 205.225 ;
        RECT 92.130 203.280 93.500 205.170 ;
        RECT 92.130 203.225 92.360 203.280 ;
        RECT 93.270 203.225 93.500 203.280 ;
        RECT 93.710 205.170 93.940 205.225 ;
        RECT 94.080 205.170 94.360 207.430 ;
        RECT 95.380 207.370 95.610 207.430 ;
        RECT 95.820 208.310 96.050 208.370 ;
        RECT 96.960 208.310 97.190 208.370 ;
        RECT 95.820 207.430 96.460 208.310 ;
        RECT 95.820 207.370 96.050 207.430 ;
        RECT 95.570 207.200 95.860 207.210 ;
        RECT 95.550 205.440 95.880 207.200 ;
        RECT 96.200 206.500 96.460 207.430 ;
        RECT 96.640 207.430 97.190 208.310 ;
        RECT 96.170 206.150 96.500 206.500 ;
        RECT 95.570 205.430 95.860 205.440 ;
        RECT 95.380 205.170 95.610 205.225 ;
        RECT 93.710 203.280 94.360 205.170 ;
        RECT 94.820 203.280 95.610 205.170 ;
        RECT 93.710 203.225 93.940 203.280 ;
        RECT 90.280 202.740 92.190 203.020 ;
        RECT 93.460 203.010 93.750 203.020 ;
        RECT 93.440 202.740 93.770 203.010 ;
        RECT 94.820 202.530 95.150 203.280 ;
        RECT 95.380 203.225 95.610 203.280 ;
        RECT 95.820 205.160 96.050 205.225 ;
        RECT 96.200 205.160 96.460 206.150 ;
        RECT 95.820 203.280 96.460 205.160 ;
        RECT 96.640 205.160 96.820 207.430 ;
        RECT 96.960 207.370 97.190 207.430 ;
        RECT 97.400 208.310 97.630 208.370 ;
        RECT 98.540 208.310 98.770 208.370 ;
        RECT 97.400 207.430 98.770 208.310 ;
        RECT 97.400 207.370 97.630 207.430 ;
        RECT 97.130 206.160 97.460 207.210 ;
        RECT 97.130 205.430 97.460 205.710 ;
        RECT 96.960 205.160 97.190 205.225 ;
        RECT 96.640 203.280 97.190 205.160 ;
        RECT 95.820 203.225 96.050 203.280 ;
        RECT 96.960 203.225 97.190 203.280 ;
        RECT 97.400 205.170 97.630 205.225 ;
        RECT 97.770 205.170 98.400 207.430 ;
        RECT 98.540 207.370 98.770 207.430 ;
        RECT 98.980 208.310 99.210 208.370 ;
        RECT 100.130 208.320 100.430 209.020 ;
        RECT 100.830 208.520 101.130 208.820 ;
        RECT 100.650 208.320 100.880 208.370 ;
        RECT 98.980 207.430 99.630 208.310 ;
        RECT 98.980 207.370 99.210 207.430 ;
        RECT 98.730 207.190 99.020 207.210 ;
        RECT 98.710 206.930 99.040 207.190 ;
        RECT 98.710 205.430 99.040 206.480 ;
        RECT 98.540 205.170 98.770 205.225 ;
        RECT 97.400 203.280 98.770 205.170 ;
        RECT 97.400 203.225 97.630 203.280 ;
        RECT 98.540 203.225 98.770 203.280 ;
        RECT 98.980 205.170 99.210 205.225 ;
        RECT 99.350 205.170 99.630 207.430 ;
        RECT 100.130 207.420 100.880 208.320 ;
        RECT 100.650 207.370 100.880 207.420 ;
        RECT 101.090 208.320 101.320 208.370 ;
        RECT 102.230 208.320 102.530 209.020 ;
        RECT 102.930 208.520 103.230 208.820 ;
        RECT 102.750 208.320 102.980 208.370 ;
        RECT 101.090 207.420 101.730 208.320 ;
        RECT 102.230 207.420 102.980 208.320 ;
        RECT 101.090 207.370 101.320 207.420 ;
        RECT 100.830 206.520 101.130 207.220 ;
        RECT 100.130 206.120 101.130 206.520 ;
        RECT 100.830 205.420 101.130 206.120 ;
        RECT 101.530 206.520 101.730 207.420 ;
        RECT 102.750 207.370 102.980 207.420 ;
        RECT 103.190 208.320 103.420 208.370 ;
        RECT 103.190 207.420 103.830 208.320 ;
        RECT 103.190 207.370 103.420 207.420 ;
        RECT 102.930 206.520 103.230 207.220 ;
        RECT 101.530 206.120 103.230 206.520 ;
        RECT 100.650 205.220 100.880 205.225 ;
        RECT 98.980 203.280 99.630 205.170 ;
        RECT 100.130 203.320 100.880 205.220 ;
        RECT 98.980 203.225 99.210 203.280 ;
        RECT 95.550 202.740 97.460 203.020 ;
        RECT 98.730 203.010 99.020 203.020 ;
        RECT 98.710 202.740 99.040 203.010 ;
        RECT 100.130 202.530 100.430 203.320 ;
        RECT 100.650 203.225 100.880 203.320 ;
        RECT 101.090 205.220 101.320 205.225 ;
        RECT 101.530 205.220 101.730 206.120 ;
        RECT 102.930 205.420 103.230 206.120 ;
        RECT 103.630 206.520 103.830 207.420 ;
        RECT 105.610 206.520 106.080 207.320 ;
        RECT 103.630 206.120 106.080 206.520 ;
        RECT 102.750 205.220 102.980 205.225 ;
        RECT 101.090 203.320 101.730 205.220 ;
        RECT 102.230 203.320 102.980 205.220 ;
        RECT 101.090 203.225 101.320 203.320 ;
        RECT 100.830 202.720 101.130 203.020 ;
        RECT 102.230 202.530 102.530 203.320 ;
        RECT 102.750 203.225 102.980 203.320 ;
        RECT 103.190 205.220 103.420 205.225 ;
        RECT 103.630 205.220 103.830 206.120 ;
        RECT 103.190 203.320 103.830 205.220 ;
        RECT 103.190 203.225 103.420 203.320 ;
        RECT 102.930 202.720 103.230 203.020 ;
        RECT 67.410 201.980 78.940 202.240 ;
        RECT 67.410 201.690 67.770 201.980 ;
        RECT 73.020 201.690 74.390 201.980 ;
        RECT 59.200 201.630 59.430 201.690 ;
        RECT 60.500 201.630 60.730 201.690 ;
        RECT 66.050 201.630 66.280 201.690 ;
        RECT 67.470 201.630 67.700 201.690 ;
        RECT 73.020 201.630 73.250 201.690 ;
        RECT 74.160 201.630 74.390 201.690 ;
        RECT 78.710 201.630 78.940 201.980 ;
        RECT 85.180 201.730 104.140 202.530 ;
        RECT 28.120 201.350 32.120 201.580 ;
        RECT 33.970 201.350 38.970 201.580 ;
        RECT 40.940 201.350 45.940 201.580 ;
        RECT 47.630 201.350 51.630 201.580 ;
        RECT 55.040 201.350 59.040 201.580 ;
        RECT 60.890 201.350 65.890 201.580 ;
        RECT 67.860 201.350 72.860 201.580 ;
        RECT 74.550 201.350 78.550 201.580 ;
        RECT 28.430 200.980 31.800 201.350 ;
        RECT 34.720 200.980 38.090 201.350 ;
        RECT 41.830 200.980 45.200 201.350 ;
        RECT 55.350 200.980 58.720 201.350 ;
        RECT 61.640 200.980 65.010 201.350 ;
        RECT 68.750 200.980 72.120 201.350 ;
        RECT 27.070 200.810 79.600 200.980 ;
        RECT 27.070 198.580 32.990 200.810 ;
        RECT 33.980 200.440 38.960 200.460 ;
        RECT 40.950 200.440 45.930 200.460 ;
        RECT 33.970 200.210 38.970 200.440 ;
        RECT 40.940 200.210 45.940 200.440 ;
        RECT 33.980 200.200 38.960 200.210 ;
        RECT 40.950 200.200 45.930 200.210 ;
        RECT 33.580 199.820 33.810 200.160 ;
        RECT 39.130 200.100 39.360 200.160 ;
        RECT 40.550 200.100 40.780 200.160 ;
        RECT 39.060 199.820 39.420 200.100 ;
        RECT 33.580 199.560 39.420 199.820 ;
        RECT 33.580 199.200 33.810 199.560 ;
        RECT 39.060 199.260 39.420 199.560 ;
        RECT 40.490 199.820 40.850 200.100 ;
        RECT 46.100 199.820 46.330 200.160 ;
        RECT 40.490 199.560 46.330 199.820 ;
        RECT 40.490 199.260 40.850 199.560 ;
        RECT 39.130 199.200 39.360 199.260 ;
        RECT 40.550 199.200 40.780 199.260 ;
        RECT 46.100 199.200 46.330 199.560 ;
        RECT 33.970 198.920 38.970 199.150 ;
        RECT 40.940 198.920 45.940 199.150 ;
        RECT 34.030 198.580 38.910 198.920 ;
        RECT 41.000 198.580 45.880 198.920 ;
        RECT 46.760 198.580 59.910 200.810 ;
        RECT 60.900 200.440 65.880 200.460 ;
        RECT 67.870 200.440 72.850 200.460 ;
        RECT 60.890 200.210 65.890 200.440 ;
        RECT 67.860 200.210 72.860 200.440 ;
        RECT 60.900 200.200 65.880 200.210 ;
        RECT 67.870 200.200 72.850 200.210 ;
        RECT 60.500 199.820 60.730 200.160 ;
        RECT 66.050 200.100 66.280 200.160 ;
        RECT 67.470 200.100 67.700 200.160 ;
        RECT 65.980 199.820 66.340 200.100 ;
        RECT 60.500 199.560 66.340 199.820 ;
        RECT 60.500 199.200 60.730 199.560 ;
        RECT 65.980 199.260 66.340 199.560 ;
        RECT 67.410 199.820 67.770 200.100 ;
        RECT 73.020 199.820 73.250 200.160 ;
        RECT 67.410 199.560 73.250 199.820 ;
        RECT 67.410 199.260 67.770 199.560 ;
        RECT 66.050 199.200 66.280 199.260 ;
        RECT 67.470 199.200 67.700 199.260 ;
        RECT 73.020 199.200 73.250 199.560 ;
        RECT 60.890 198.920 65.890 199.150 ;
        RECT 67.860 198.920 72.860 199.150 ;
        RECT 60.950 198.580 65.830 198.920 ;
        RECT 67.920 198.580 72.800 198.920 ;
        RECT 73.680 198.580 79.600 200.810 ;
        RECT 85.380 200.940 85.680 201.730 ;
        RECT 86.080 201.240 86.380 201.540 ;
        RECT 85.900 200.940 86.130 201.035 ;
        RECT 85.380 199.040 86.130 200.940 ;
        RECT 85.900 199.035 86.130 199.040 ;
        RECT 86.340 200.940 86.570 201.035 ;
        RECT 87.480 200.940 87.780 201.730 ;
        RECT 88.180 201.240 88.480 201.540 ;
        RECT 88.000 200.940 88.230 201.035 ;
        RECT 86.340 199.040 86.980 200.940 ;
        RECT 87.480 199.040 88.230 200.940 ;
        RECT 86.340 199.035 86.570 199.040 ;
        RECT 27.070 197.820 79.600 198.580 ;
        RECT 24.010 195.300 25.830 197.310 ;
        RECT 27.070 195.590 32.990 197.820 ;
        RECT 34.030 197.480 38.910 197.820 ;
        RECT 41.000 197.480 45.880 197.820 ;
        RECT 33.970 197.250 38.970 197.480 ;
        RECT 40.940 197.250 45.940 197.480 ;
        RECT 33.580 196.840 33.810 197.200 ;
        RECT 39.130 197.140 39.360 197.200 ;
        RECT 40.550 197.140 40.780 197.200 ;
        RECT 39.060 196.840 39.420 197.140 ;
        RECT 33.580 196.580 39.420 196.840 ;
        RECT 33.580 196.240 33.810 196.580 ;
        RECT 39.060 196.300 39.420 196.580 ;
        RECT 40.490 196.840 40.850 197.140 ;
        RECT 46.100 196.840 46.330 197.200 ;
        RECT 40.490 196.580 46.330 196.840 ;
        RECT 40.490 196.300 40.850 196.580 ;
        RECT 39.130 196.240 39.360 196.300 ;
        RECT 40.550 196.240 40.780 196.300 ;
        RECT 46.100 196.240 46.330 196.580 ;
        RECT 33.980 196.190 38.960 196.200 ;
        RECT 40.950 196.190 45.930 196.200 ;
        RECT 33.970 195.960 38.970 196.190 ;
        RECT 40.940 195.960 45.940 196.190 ;
        RECT 33.980 195.940 38.960 195.960 ;
        RECT 40.950 195.940 45.930 195.960 ;
        RECT 46.760 195.590 59.910 197.820 ;
        RECT 60.950 197.480 65.830 197.820 ;
        RECT 67.920 197.480 72.800 197.820 ;
        RECT 60.890 197.250 65.890 197.480 ;
        RECT 67.860 197.250 72.860 197.480 ;
        RECT 60.500 196.840 60.730 197.200 ;
        RECT 66.050 197.140 66.280 197.200 ;
        RECT 67.470 197.140 67.700 197.200 ;
        RECT 65.980 196.840 66.340 197.140 ;
        RECT 60.500 196.580 66.340 196.840 ;
        RECT 60.500 196.240 60.730 196.580 ;
        RECT 65.980 196.300 66.340 196.580 ;
        RECT 67.410 196.840 67.770 197.140 ;
        RECT 73.020 196.840 73.250 197.200 ;
        RECT 67.410 196.580 73.250 196.840 ;
        RECT 67.410 196.300 67.770 196.580 ;
        RECT 66.050 196.240 66.280 196.300 ;
        RECT 67.470 196.240 67.700 196.300 ;
        RECT 73.020 196.240 73.250 196.580 ;
        RECT 60.900 196.190 65.880 196.200 ;
        RECT 67.870 196.190 72.850 196.200 ;
        RECT 60.890 195.960 65.890 196.190 ;
        RECT 67.860 195.960 72.860 196.190 ;
        RECT 60.900 195.940 65.880 195.960 ;
        RECT 67.870 195.940 72.850 195.960 ;
        RECT 73.680 195.590 79.600 197.820 ;
        RECT 83.350 198.140 85.410 198.380 ;
        RECT 86.080 198.140 86.380 198.840 ;
        RECT 83.350 197.740 86.380 198.140 ;
        RECT 83.350 197.610 85.410 197.740 ;
        RECT 83.350 197.600 84.940 197.610 ;
        RECT 86.080 197.040 86.380 197.740 ;
        RECT 86.780 198.140 86.980 199.040 ;
        RECT 88.000 199.035 88.230 199.040 ;
        RECT 88.440 200.940 88.670 201.035 ;
        RECT 89.550 200.980 89.880 201.730 ;
        RECT 90.280 201.240 92.190 201.520 ;
        RECT 93.440 201.250 93.770 201.520 ;
        RECT 93.460 201.240 93.750 201.250 ;
        RECT 90.110 200.980 90.340 201.035 ;
        RECT 88.440 199.040 89.080 200.940 ;
        RECT 89.550 199.090 90.340 200.980 ;
        RECT 88.440 199.035 88.670 199.040 ;
        RECT 88.180 198.140 88.480 198.840 ;
        RECT 86.780 197.740 88.480 198.140 ;
        RECT 85.900 196.840 86.130 196.890 ;
        RECT 27.070 195.420 79.600 195.590 ;
        RECT 85.380 195.940 86.130 196.840 ;
        RECT 28.430 195.050 31.800 195.420 ;
        RECT 34.720 195.050 38.090 195.420 ;
        RECT 41.830 195.050 45.200 195.420 ;
        RECT 55.350 195.050 58.720 195.420 ;
        RECT 61.640 195.050 65.010 195.420 ;
        RECT 68.750 195.050 72.120 195.420 ;
        RECT 85.380 195.240 85.680 195.940 ;
        RECT 85.900 195.890 86.130 195.940 ;
        RECT 86.340 196.840 86.570 196.890 ;
        RECT 86.780 196.840 86.980 197.740 ;
        RECT 88.180 197.040 88.480 197.740 ;
        RECT 88.880 198.140 89.080 199.040 ;
        RECT 90.110 199.035 90.340 199.090 ;
        RECT 90.550 200.980 90.780 201.035 ;
        RECT 91.690 200.980 91.920 201.035 ;
        RECT 90.550 199.100 91.190 200.980 ;
        RECT 90.550 199.035 90.780 199.100 ;
        RECT 90.300 198.820 90.590 198.830 ;
        RECT 88.880 197.740 89.280 198.140 ;
        RECT 88.000 196.840 88.230 196.890 ;
        RECT 86.340 195.940 86.980 196.840 ;
        RECT 87.480 195.940 88.230 196.840 ;
        RECT 86.340 195.890 86.570 195.940 ;
        RECT 86.080 195.440 86.380 195.740 ;
        RECT 87.480 195.240 87.780 195.940 ;
        RECT 88.000 195.890 88.230 195.940 ;
        RECT 88.440 196.840 88.670 196.890 ;
        RECT 88.880 196.840 89.080 197.740 ;
        RECT 90.280 197.060 90.610 198.820 ;
        RECT 90.930 198.110 91.190 199.100 ;
        RECT 91.370 199.100 91.920 200.980 ;
        RECT 90.900 197.760 91.230 198.110 ;
        RECT 90.300 197.050 90.590 197.060 ;
        RECT 88.440 195.940 89.080 196.840 ;
        RECT 90.110 196.830 90.340 196.890 ;
        RECT 89.520 195.950 90.340 196.830 ;
        RECT 88.440 195.890 88.670 195.940 ;
        RECT 88.180 195.440 88.480 195.740 ;
        RECT 89.520 195.240 89.810 195.950 ;
        RECT 90.110 195.890 90.340 195.950 ;
        RECT 90.550 196.830 90.780 196.890 ;
        RECT 90.930 196.830 91.190 197.760 ;
        RECT 90.550 195.950 91.190 196.830 ;
        RECT 91.370 196.830 91.550 199.100 ;
        RECT 91.690 199.035 91.920 199.100 ;
        RECT 92.130 200.980 92.360 201.035 ;
        RECT 93.270 200.980 93.500 201.035 ;
        RECT 92.130 199.090 93.500 200.980 ;
        RECT 92.130 199.035 92.360 199.090 ;
        RECT 91.860 198.550 92.190 198.830 ;
        RECT 91.860 197.050 92.190 198.100 ;
        RECT 91.690 196.830 91.920 196.890 ;
        RECT 91.370 195.950 91.920 196.830 ;
        RECT 90.550 195.890 90.780 195.950 ;
        RECT 91.690 195.890 91.920 195.950 ;
        RECT 92.130 196.830 92.360 196.890 ;
        RECT 92.500 196.830 93.130 199.090 ;
        RECT 93.270 199.035 93.500 199.090 ;
        RECT 93.710 200.980 93.940 201.035 ;
        RECT 93.710 199.090 94.360 200.980 ;
        RECT 93.710 199.035 93.940 199.090 ;
        RECT 93.440 197.780 93.770 198.830 ;
        RECT 93.440 197.070 93.770 197.330 ;
        RECT 93.460 197.050 93.750 197.070 ;
        RECT 93.270 196.830 93.500 196.890 ;
        RECT 92.130 195.950 93.500 196.830 ;
        RECT 92.130 195.890 92.360 195.950 ;
        RECT 93.270 195.890 93.500 195.950 ;
        RECT 93.710 196.830 93.940 196.890 ;
        RECT 94.080 196.830 94.360 199.090 ;
        RECT 100.130 200.940 100.430 201.730 ;
        RECT 100.830 201.240 101.130 201.540 ;
        RECT 100.650 200.940 100.880 201.035 ;
        RECT 100.130 199.040 100.880 200.940 ;
        RECT 100.650 199.035 100.880 199.040 ;
        RECT 101.090 200.940 101.320 201.035 ;
        RECT 102.230 200.940 102.530 201.730 ;
        RECT 102.930 201.240 103.230 201.540 ;
        RECT 102.750 200.940 102.980 201.035 ;
        RECT 101.090 199.040 101.730 200.940 ;
        RECT 102.230 199.040 102.980 200.940 ;
        RECT 101.090 199.035 101.320 199.040 ;
        RECT 98.720 198.140 99.400 198.220 ;
        RECT 100.830 198.140 101.130 198.840 ;
        RECT 98.720 197.740 101.130 198.140 ;
        RECT 98.720 197.280 99.400 197.740 ;
        RECT 100.830 197.040 101.130 197.740 ;
        RECT 101.530 198.140 101.730 199.040 ;
        RECT 102.750 199.035 102.980 199.040 ;
        RECT 103.190 200.940 103.420 201.035 ;
        RECT 103.190 199.040 103.830 200.940 ;
        RECT 103.190 199.035 103.420 199.040 ;
        RECT 102.930 198.140 103.230 198.840 ;
        RECT 101.530 197.740 103.230 198.140 ;
        RECT 100.650 196.840 100.880 196.890 ;
        RECT 93.710 195.950 94.360 196.830 ;
        RECT 93.710 195.890 93.940 195.950 ;
        RECT 100.130 195.940 100.880 196.840 ;
        RECT 90.300 195.720 90.590 195.730 ;
        RECT 91.880 195.720 92.170 195.730 ;
        RECT 93.460 195.720 93.750 195.730 ;
        RECT 90.180 195.390 90.710 195.720 ;
        RECT 91.860 195.450 92.190 195.720 ;
        RECT 93.330 195.390 93.860 195.720 ;
        RECT 100.130 195.240 100.430 195.940 ;
        RECT 100.650 195.890 100.880 195.940 ;
        RECT 101.090 196.840 101.320 196.890 ;
        RECT 101.530 196.840 101.730 197.740 ;
        RECT 102.930 197.040 103.230 197.740 ;
        RECT 103.630 198.140 103.830 199.040 ;
        RECT 107.100 198.140 107.570 198.930 ;
        RECT 103.630 197.740 107.570 198.140 ;
        RECT 102.750 196.840 102.980 196.890 ;
        RECT 101.090 195.940 101.730 196.840 ;
        RECT 102.230 195.940 102.980 196.840 ;
        RECT 101.090 195.890 101.320 195.940 ;
        RECT 100.830 195.440 101.130 195.740 ;
        RECT 102.230 195.240 102.530 195.940 ;
        RECT 102.750 195.890 102.980 195.940 ;
        RECT 103.190 196.840 103.420 196.890 ;
        RECT 103.630 196.840 103.830 197.740 ;
        RECT 103.190 195.940 103.830 196.840 ;
        RECT 103.190 195.890 103.420 195.940 ;
        RECT 102.930 195.440 103.230 195.740 ;
        RECT 28.120 194.820 32.120 195.050 ;
        RECT 33.970 194.820 38.970 195.050 ;
        RECT 40.940 194.820 45.940 195.050 ;
        RECT 47.630 194.820 51.630 195.050 ;
        RECT 55.040 194.820 59.040 195.050 ;
        RECT 60.890 194.820 65.890 195.050 ;
        RECT 67.860 194.820 72.860 195.050 ;
        RECT 74.550 194.820 78.550 195.050 ;
        RECT 27.730 194.420 27.960 194.770 ;
        RECT 32.280 194.710 32.510 194.770 ;
        RECT 33.580 194.710 33.810 194.770 ;
        RECT 39.130 194.710 39.360 194.770 ;
        RECT 40.550 194.710 40.780 194.770 ;
        RECT 46.100 194.710 46.330 194.770 ;
        RECT 47.240 194.710 47.470 194.770 ;
        RECT 32.280 194.420 33.810 194.710 ;
        RECT 39.060 194.420 39.420 194.710 ;
        RECT 27.730 194.160 39.420 194.420 ;
        RECT 27.730 193.770 27.960 194.160 ;
        RECT 32.280 193.870 33.810 194.160 ;
        RECT 39.060 193.870 39.420 194.160 ;
        RECT 40.490 194.420 40.850 194.710 ;
        RECT 46.100 194.420 47.470 194.710 ;
        RECT 51.790 194.420 52.020 194.770 ;
        RECT 40.490 194.160 52.020 194.420 ;
        RECT 40.490 193.870 40.850 194.160 ;
        RECT 46.100 193.870 47.470 194.160 ;
        RECT 32.280 193.770 32.510 193.870 ;
        RECT 33.580 193.810 33.810 193.870 ;
        RECT 39.130 193.810 39.360 193.870 ;
        RECT 40.550 193.810 40.780 193.870 ;
        RECT 46.100 193.810 46.330 193.870 ;
        RECT 47.240 193.810 47.470 193.870 ;
        RECT 47.270 193.790 47.470 193.810 ;
        RECT 47.270 193.770 47.630 193.790 ;
        RECT 51.790 193.770 52.020 194.160 ;
        RECT 27.730 193.530 32.510 193.770 ;
        RECT 33.980 193.760 38.960 193.770 ;
        RECT 40.950 193.760 45.930 193.770 ;
        RECT 33.970 193.530 38.970 193.760 ;
        RECT 40.940 193.530 45.940 193.760 ;
        RECT 27.730 193.510 32.110 193.530 ;
        RECT 33.980 193.510 38.960 193.530 ;
        RECT 40.950 193.510 45.930 193.530 ;
        RECT 47.270 193.510 52.020 193.770 ;
        RECT 54.650 194.420 54.880 194.770 ;
        RECT 59.200 194.710 59.430 194.770 ;
        RECT 60.500 194.710 60.730 194.770 ;
        RECT 66.050 194.710 66.280 194.770 ;
        RECT 67.470 194.710 67.700 194.770 ;
        RECT 73.020 194.710 73.250 194.770 ;
        RECT 74.160 194.710 74.390 194.770 ;
        RECT 59.200 194.420 60.730 194.710 ;
        RECT 65.980 194.420 66.340 194.710 ;
        RECT 54.650 194.160 66.340 194.420 ;
        RECT 54.650 193.770 54.880 194.160 ;
        RECT 59.200 193.870 60.730 194.160 ;
        RECT 65.980 193.870 66.340 194.160 ;
        RECT 67.410 194.420 67.770 194.710 ;
        RECT 73.020 194.420 74.390 194.710 ;
        RECT 78.710 194.420 78.940 194.770 ;
        RECT 85.180 194.440 104.140 195.240 ;
        RECT 67.410 194.160 78.940 194.420 ;
        RECT 67.410 193.870 67.770 194.160 ;
        RECT 73.020 193.870 74.390 194.160 ;
        RECT 59.200 193.770 59.430 193.870 ;
        RECT 60.500 193.810 60.730 193.870 ;
        RECT 66.050 193.810 66.280 193.870 ;
        RECT 67.470 193.810 67.700 193.870 ;
        RECT 73.020 193.810 73.250 193.870 ;
        RECT 74.160 193.810 74.390 193.870 ;
        RECT 74.190 193.790 74.390 193.810 ;
        RECT 74.190 193.770 74.550 193.790 ;
        RECT 78.710 193.770 78.940 194.160 ;
        RECT 54.650 193.530 59.430 193.770 ;
        RECT 60.900 193.760 65.880 193.770 ;
        RECT 67.870 193.760 72.850 193.770 ;
        RECT 60.890 193.530 65.890 193.760 ;
        RECT 67.860 193.530 72.860 193.760 ;
        RECT 54.650 193.510 59.030 193.530 ;
        RECT 60.900 193.510 65.880 193.530 ;
        RECT 67.870 193.510 72.850 193.530 ;
        RECT 74.190 193.510 78.940 193.770 ;
        RECT 85.380 193.740 85.680 194.440 ;
        RECT 86.080 193.940 86.380 194.240 ;
        RECT 85.900 193.740 86.130 193.790 ;
        RECT 85.380 192.840 86.130 193.740 ;
        RECT 29.210 192.390 49.330 192.650 ;
        RECT 20.500 191.850 22.660 192.070 ;
        RECT 30.410 191.990 50.530 192.250 ;
        RECT 53.000 191.850 53.640 192.820 ;
        RECT 85.900 192.790 86.130 192.840 ;
        RECT 86.340 193.740 86.570 193.790 ;
        RECT 87.480 193.740 87.780 194.440 ;
        RECT 88.180 193.940 88.480 194.240 ;
        RECT 88.000 193.740 88.230 193.790 ;
        RECT 86.340 192.840 86.980 193.740 ;
        RECT 87.480 192.840 88.230 193.740 ;
        RECT 86.340 192.790 86.570 192.840 ;
        RECT 56.130 192.390 76.250 192.650 ;
        RECT 57.330 191.990 77.450 192.250 ;
        RECT 79.210 191.940 79.980 192.100 ;
        RECT 82.410 191.940 83.520 192.260 ;
        RECT 86.080 191.940 86.380 192.640 ;
        RECT 20.500 191.590 51.040 191.850 ;
        RECT 53.000 191.590 77.960 191.850 ;
        RECT 12.770 172.620 14.930 185.210 ;
        RECT 20.500 179.480 22.660 191.590 ;
        RECT 28.390 189.480 28.580 191.590 ;
        RECT 30.420 191.020 31.140 191.070 ;
        RECT 48.610 191.020 49.330 191.040 ;
        RECT 29.195 190.790 39.190 191.020 ;
        RECT 40.555 190.790 50.550 191.020 ;
        RECT 30.420 190.760 31.140 190.790 ;
        RECT 48.610 190.780 49.330 190.790 ;
        RECT 28.720 190.430 29.040 190.740 ;
        RECT 38.480 190.380 39.200 190.430 ;
        RECT 39.340 190.410 39.680 190.760 ;
        RECT 40.070 190.410 40.410 190.760 ;
        RECT 40.560 190.380 41.280 190.430 ;
        RECT 50.710 190.400 51.040 190.760 ;
        RECT 53.000 190.440 53.640 191.590 ;
        RECT 29.195 190.150 39.200 190.380 ;
        RECT 40.555 190.150 50.550 190.380 ;
        RECT 38.480 190.110 39.200 190.150 ;
        RECT 40.560 190.100 41.280 190.150 ;
        RECT 29.220 189.820 29.940 189.870 ;
        RECT 40.550 189.820 41.610 189.840 ;
        RECT 49.810 189.820 50.530 189.880 ;
        RECT 29.195 189.590 39.190 189.820 ;
        RECT 40.550 189.590 50.550 189.820 ;
        RECT 29.220 189.550 29.940 189.590 ;
        RECT 40.550 189.580 41.610 189.590 ;
        RECT 49.810 189.540 50.530 189.590 ;
        RECT 28.740 189.480 29.020 189.540 ;
        RECT 28.390 189.290 29.020 189.480 ;
        RECT 28.390 187.080 28.580 189.290 ;
        RECT 28.740 189.230 29.020 189.290 ;
        RECT 39.380 189.230 39.650 189.540 ;
        RECT 40.100 189.230 40.380 189.540 ;
        RECT 50.740 189.480 51.010 189.540 ;
        RECT 55.310 189.480 55.500 191.590 ;
        RECT 79.210 191.540 86.380 191.940 ;
        RECT 79.210 191.410 79.980 191.540 ;
        RECT 82.410 191.240 83.520 191.540 ;
        RECT 57.340 191.020 58.060 191.070 ;
        RECT 75.530 191.020 76.250 191.040 ;
        RECT 56.115 190.790 66.110 191.020 ;
        RECT 67.475 190.790 77.470 191.020 ;
        RECT 86.080 190.840 86.380 191.540 ;
        RECT 86.780 191.940 86.980 192.840 ;
        RECT 88.000 192.790 88.230 192.840 ;
        RECT 88.440 193.740 88.670 193.790 ;
        RECT 88.440 192.840 89.080 193.740 ;
        RECT 89.970 193.235 90.970 194.190 ;
        RECT 88.440 192.790 88.670 192.840 ;
        RECT 88.180 191.940 88.480 192.640 ;
        RECT 86.780 191.540 88.480 191.940 ;
        RECT 57.340 190.760 58.060 190.790 ;
        RECT 75.530 190.780 76.250 190.790 ;
        RECT 55.640 190.430 55.960 190.740 ;
        RECT 65.400 190.380 66.120 190.430 ;
        RECT 66.260 190.410 66.600 190.760 ;
        RECT 66.990 190.410 67.330 190.760 ;
        RECT 67.480 190.380 68.200 190.430 ;
        RECT 77.630 190.400 77.960 190.760 ;
        RECT 85.900 190.640 86.130 190.645 ;
        RECT 56.115 190.150 66.120 190.380 ;
        RECT 67.475 190.150 77.470 190.380 ;
        RECT 65.400 190.110 66.120 190.150 ;
        RECT 67.480 190.100 68.200 190.150 ;
        RECT 56.140 189.820 56.860 189.870 ;
        RECT 67.470 189.820 68.530 189.840 ;
        RECT 76.730 189.820 77.450 189.880 ;
        RECT 56.115 189.590 66.110 189.820 ;
        RECT 67.470 189.590 77.470 189.820 ;
        RECT 56.140 189.550 56.860 189.590 ;
        RECT 67.470 189.580 68.530 189.590 ;
        RECT 76.730 189.540 77.450 189.590 ;
        RECT 55.660 189.480 55.940 189.540 ;
        RECT 50.740 189.290 51.370 189.480 ;
        RECT 50.740 189.230 51.010 189.290 ;
        RECT 38.480 189.180 39.200 189.230 ;
        RECT 40.560 189.180 41.610 189.210 ;
        RECT 29.195 188.950 39.200 189.180 ;
        RECT 40.555 188.950 50.550 189.180 ;
        RECT 38.480 188.910 39.200 188.950 ;
        RECT 40.560 188.900 41.280 188.950 ;
        RECT 30.420 188.620 31.140 188.670 ;
        RECT 48.610 188.620 49.330 188.640 ;
        RECT 29.195 188.390 39.190 188.620 ;
        RECT 40.555 188.390 50.550 188.620 ;
        RECT 30.420 188.360 31.140 188.390 ;
        RECT 48.610 188.380 49.330 188.390 ;
        RECT 28.720 188.030 29.040 188.340 ;
        RECT 38.480 187.980 39.200 188.030 ;
        RECT 39.340 188.010 39.680 188.360 ;
        RECT 40.070 188.010 40.410 188.360 ;
        RECT 40.560 187.980 41.280 188.030 ;
        RECT 50.710 188.000 51.040 188.360 ;
        RECT 29.195 187.750 39.200 187.980 ;
        RECT 40.555 187.750 50.550 187.980 ;
        RECT 38.480 187.710 39.200 187.750 ;
        RECT 40.560 187.700 41.280 187.750 ;
        RECT 29.220 187.420 29.940 187.470 ;
        RECT 40.550 187.420 41.650 187.440 ;
        RECT 49.810 187.420 50.530 187.480 ;
        RECT 29.195 187.190 39.190 187.420 ;
        RECT 40.550 187.190 50.550 187.420 ;
        RECT 29.220 187.150 29.940 187.190 ;
        RECT 40.550 187.180 41.650 187.190 ;
        RECT 49.810 187.140 50.530 187.190 ;
        RECT 28.740 187.080 29.020 187.140 ;
        RECT 28.390 186.890 29.020 187.080 ;
        RECT 28.740 186.830 29.020 186.890 ;
        RECT 39.380 186.830 39.650 187.140 ;
        RECT 40.100 186.830 40.380 187.140 ;
        RECT 50.740 187.080 51.010 187.140 ;
        RECT 51.180 187.080 51.370 189.290 ;
        RECT 50.740 186.890 51.370 187.080 ;
        RECT 55.310 189.290 55.940 189.480 ;
        RECT 55.310 187.080 55.500 189.290 ;
        RECT 55.660 189.230 55.940 189.290 ;
        RECT 66.300 189.230 66.570 189.540 ;
        RECT 67.020 189.230 67.300 189.540 ;
        RECT 77.660 189.480 77.930 189.540 ;
        RECT 77.660 189.290 78.290 189.480 ;
        RECT 77.660 189.230 77.930 189.290 ;
        RECT 65.400 189.180 66.120 189.230 ;
        RECT 67.480 189.180 68.530 189.210 ;
        RECT 56.115 188.950 66.120 189.180 ;
        RECT 67.475 188.950 77.470 189.180 ;
        RECT 65.400 188.910 66.120 188.950 ;
        RECT 67.480 188.900 68.200 188.950 ;
        RECT 57.340 188.620 58.060 188.670 ;
        RECT 75.530 188.620 76.250 188.640 ;
        RECT 56.115 188.390 66.110 188.620 ;
        RECT 67.475 188.390 77.470 188.620 ;
        RECT 57.340 188.360 58.060 188.390 ;
        RECT 75.530 188.380 76.250 188.390 ;
        RECT 55.640 188.030 55.960 188.340 ;
        RECT 65.400 187.980 66.120 188.030 ;
        RECT 66.260 188.010 66.600 188.360 ;
        RECT 66.990 188.010 67.330 188.360 ;
        RECT 67.480 187.980 68.200 188.030 ;
        RECT 77.630 188.000 77.960 188.360 ;
        RECT 56.115 187.750 66.120 187.980 ;
        RECT 67.475 187.750 77.470 187.980 ;
        RECT 65.400 187.710 66.120 187.750 ;
        RECT 67.480 187.700 68.200 187.750 ;
        RECT 56.140 187.420 56.860 187.470 ;
        RECT 67.470 187.420 68.570 187.440 ;
        RECT 76.730 187.420 77.450 187.480 ;
        RECT 56.115 187.190 66.110 187.420 ;
        RECT 67.470 187.190 77.470 187.420 ;
        RECT 56.140 187.150 56.860 187.190 ;
        RECT 67.470 187.180 68.570 187.190 ;
        RECT 76.730 187.140 77.450 187.190 ;
        RECT 55.660 187.080 55.940 187.140 ;
        RECT 55.310 186.890 55.940 187.080 ;
        RECT 50.740 186.830 51.010 186.890 ;
        RECT 38.480 186.780 39.200 186.830 ;
        RECT 40.560 186.780 41.650 186.810 ;
        RECT 24.490 185.900 25.220 186.650 ;
        RECT 29.195 186.550 39.200 186.780 ;
        RECT 40.555 186.550 50.550 186.780 ;
        RECT 38.480 186.510 39.200 186.550 ;
        RECT 40.560 186.540 41.260 186.550 ;
        RECT 51.180 185.900 51.370 186.890 ;
        RECT 55.660 186.830 55.940 186.890 ;
        RECT 66.300 186.830 66.570 187.140 ;
        RECT 67.020 186.830 67.300 187.140 ;
        RECT 77.660 187.080 77.930 187.140 ;
        RECT 78.100 187.080 78.290 189.290 ;
        RECT 85.380 188.740 86.130 190.640 ;
        RECT 85.380 187.950 85.680 188.740 ;
        RECT 85.900 188.645 86.130 188.740 ;
        RECT 86.340 190.640 86.570 190.645 ;
        RECT 86.780 190.640 86.980 191.540 ;
        RECT 88.180 190.840 88.480 191.540 ;
        RECT 88.880 191.940 89.080 192.840 ;
        RECT 89.970 191.940 90.970 192.235 ;
        RECT 88.880 191.540 90.970 191.940 ;
        RECT 88.000 190.640 88.230 190.645 ;
        RECT 86.340 188.740 86.980 190.640 ;
        RECT 87.480 188.740 88.230 190.640 ;
        RECT 86.340 188.645 86.570 188.740 ;
        RECT 86.080 188.140 86.380 188.440 ;
        RECT 87.480 187.950 87.780 188.740 ;
        RECT 88.000 188.645 88.230 188.740 ;
        RECT 88.440 190.640 88.670 190.645 ;
        RECT 88.880 190.640 89.080 191.540 ;
        RECT 88.440 188.740 89.080 190.640 ;
        RECT 88.440 188.645 88.670 188.740 ;
        RECT 88.180 188.140 88.480 188.440 ;
        RECT 85.180 187.150 104.140 187.950 ;
        RECT 77.660 186.890 78.290 187.080 ;
        RECT 77.660 186.830 77.930 186.890 ;
        RECT 65.400 186.780 66.120 186.830 ;
        RECT 67.480 186.780 68.570 186.810 ;
        RECT 56.115 186.550 66.120 186.780 ;
        RECT 67.475 186.550 77.470 186.780 ;
        RECT 65.400 186.510 66.120 186.550 ;
        RECT 67.480 186.540 68.180 186.550 ;
        RECT 78.100 185.900 78.290 186.890 ;
        RECT 24.490 185.640 51.370 185.900 ;
        RECT 53.940 185.640 78.290 185.900 ;
        RECT 85.380 186.360 85.680 187.150 ;
        RECT 86.080 186.660 86.380 186.960 ;
        RECT 85.900 186.360 86.130 186.455 ;
        RECT 24.490 184.620 25.220 185.640 ;
        RECT 53.940 185.170 54.180 185.640 ;
        RECT 51.080 184.990 54.180 185.170 ;
        RECT 34.985 184.570 44.985 184.800 ;
        RECT 34.995 184.540 44.975 184.570 ;
        RECT 34.550 184.460 34.780 184.520 ;
        RECT 45.190 184.460 45.420 184.520 ;
        RECT 34.480 183.620 34.840 184.460 ;
        RECT 45.120 183.620 45.480 184.460 ;
        RECT 34.550 183.560 34.780 183.620 ;
        RECT 45.190 183.560 45.420 183.620 ;
        RECT 34.985 183.280 44.985 183.510 ;
        RECT 51.080 183.140 51.810 184.990 ;
        RECT 61.905 184.570 71.905 184.800 ;
        RECT 61.915 184.540 71.895 184.570 ;
        RECT 61.470 184.460 61.700 184.520 ;
        RECT 72.110 184.460 72.340 184.520 ;
        RECT 85.380 184.460 86.130 186.360 ;
        RECT 61.400 183.620 61.760 184.460 ;
        RECT 72.040 183.620 72.400 184.460 ;
        RECT 85.900 184.455 86.130 184.460 ;
        RECT 86.340 186.360 86.570 186.455 ;
        RECT 87.480 186.360 87.780 187.150 ;
        RECT 88.180 186.660 88.480 186.960 ;
        RECT 88.000 186.360 88.230 186.455 ;
        RECT 86.340 184.460 86.980 186.360 ;
        RECT 87.480 184.460 88.230 186.360 ;
        RECT 86.340 184.455 86.570 184.460 ;
        RECT 61.470 183.560 61.700 183.620 ;
        RECT 72.110 183.560 72.340 183.620 ;
        RECT 81.570 183.560 83.430 183.870 ;
        RECT 86.080 183.560 86.380 184.260 ;
        RECT 61.905 183.280 71.905 183.510 ;
        RECT 81.570 183.160 86.380 183.560 ;
        RECT 81.570 182.920 83.430 183.160 ;
        RECT 27.070 182.300 79.600 182.660 ;
        RECT 86.080 182.460 86.380 183.160 ;
        RECT 86.780 183.560 86.980 184.460 ;
        RECT 88.000 184.455 88.230 184.460 ;
        RECT 88.440 186.360 88.670 186.455 ;
        RECT 88.440 184.460 89.080 186.360 ;
        RECT 88.440 184.455 88.670 184.460 ;
        RECT 88.180 183.560 88.480 184.260 ;
        RECT 86.780 183.160 88.480 183.560 ;
        RECT 27.070 180.070 30.310 182.300 ;
        RECT 30.610 181.680 39.480 181.940 ;
        RECT 40.710 181.930 48.690 181.940 ;
        RECT 40.705 181.700 48.705 181.930 ;
        RECT 40.710 181.680 48.690 181.700 ;
        RECT 30.610 181.290 30.840 181.680 ;
        RECT 39.250 181.590 39.480 181.680 ;
        RECT 40.270 181.590 40.500 181.650 ;
        RECT 39.250 181.290 40.500 181.590 ;
        RECT 48.910 181.290 49.140 181.650 ;
        RECT 30.610 181.030 49.140 181.290 ;
        RECT 30.610 180.690 30.840 181.030 ;
        RECT 39.250 180.750 40.500 181.030 ;
        RECT 39.250 180.690 39.480 180.750 ;
        RECT 40.270 180.690 40.500 180.750 ;
        RECT 48.910 180.690 49.140 181.030 ;
        RECT 31.045 180.410 39.045 180.640 ;
        RECT 40.705 180.410 48.705 180.640 ;
        RECT 31.105 180.070 38.985 180.410 ;
        RECT 40.765 180.070 48.645 180.410 ;
        RECT 49.430 180.070 57.230 182.300 ;
        RECT 57.530 181.680 66.400 181.940 ;
        RECT 67.630 181.930 75.610 181.940 ;
        RECT 67.625 181.700 75.625 181.930 ;
        RECT 67.630 181.680 75.610 181.700 ;
        RECT 57.530 181.290 57.760 181.680 ;
        RECT 66.170 181.590 66.400 181.680 ;
        RECT 67.190 181.590 67.420 181.650 ;
        RECT 66.170 181.290 67.420 181.590 ;
        RECT 75.830 181.290 76.060 181.650 ;
        RECT 57.530 181.030 76.060 181.290 ;
        RECT 57.530 180.690 57.760 181.030 ;
        RECT 66.170 180.750 67.420 181.030 ;
        RECT 66.170 180.690 66.400 180.750 ;
        RECT 67.190 180.690 67.420 180.750 ;
        RECT 75.830 180.690 76.060 181.030 ;
        RECT 57.965 180.410 65.965 180.640 ;
        RECT 67.625 180.410 75.625 180.640 ;
        RECT 58.025 180.070 65.905 180.410 ;
        RECT 67.685 180.070 75.565 180.410 ;
        RECT 76.360 180.070 79.600 182.300 ;
        RECT 85.900 182.260 86.130 182.310 ;
        RECT 85.380 181.360 86.130 182.260 ;
        RECT 85.380 180.660 85.680 181.360 ;
        RECT 85.900 181.310 86.130 181.360 ;
        RECT 86.340 182.260 86.570 182.310 ;
        RECT 86.780 182.260 86.980 183.160 ;
        RECT 88.180 182.460 88.480 183.160 ;
        RECT 88.880 183.560 89.080 184.460 ;
        RECT 88.880 183.160 89.280 183.560 ;
        RECT 88.000 182.260 88.230 182.310 ;
        RECT 86.340 181.360 86.980 182.260 ;
        RECT 87.480 181.360 88.230 182.260 ;
        RECT 86.340 181.310 86.570 181.360 ;
        RECT 86.080 180.860 86.380 181.160 ;
        RECT 87.480 180.660 87.780 181.360 ;
        RECT 88.000 181.310 88.230 181.360 ;
        RECT 88.440 182.260 88.670 182.310 ;
        RECT 88.880 182.260 89.080 183.160 ;
        RECT 88.440 181.360 89.080 182.260 ;
        RECT 88.440 181.310 88.670 181.360 ;
        RECT 88.180 180.860 88.480 181.160 ;
        RECT 27.070 179.310 79.600 180.070 ;
        RECT 85.180 179.860 104.140 180.660 ;
        RECT 12.770 158.900 14.930 171.490 ;
        RECT 20.500 167.790 22.660 178.350 ;
        RECT 27.070 177.080 30.310 179.310 ;
        RECT 31.105 178.970 38.985 179.310 ;
        RECT 40.765 178.970 48.645 179.310 ;
        RECT 31.045 178.740 39.045 178.970 ;
        RECT 40.705 178.740 48.705 178.970 ;
        RECT 30.610 178.350 30.840 178.690 ;
        RECT 39.250 178.630 39.480 178.690 ;
        RECT 40.270 178.630 40.500 178.690 ;
        RECT 39.250 178.350 40.500 178.630 ;
        RECT 48.910 178.350 49.140 178.690 ;
        RECT 30.610 178.090 49.140 178.350 ;
        RECT 30.610 177.700 30.840 178.090 ;
        RECT 39.250 177.790 40.500 178.090 ;
        RECT 39.250 177.700 39.480 177.790 ;
        RECT 40.270 177.730 40.500 177.790 ;
        RECT 48.910 177.730 49.140 178.090 ;
        RECT 30.610 177.440 39.480 177.700 ;
        RECT 40.710 177.680 48.690 177.700 ;
        RECT 40.705 177.450 48.705 177.680 ;
        RECT 40.710 177.440 48.690 177.450 ;
        RECT 49.430 177.080 57.230 179.310 ;
        RECT 58.025 178.970 65.905 179.310 ;
        RECT 67.685 178.970 75.565 179.310 ;
        RECT 57.965 178.740 65.965 178.970 ;
        RECT 67.625 178.740 75.625 178.970 ;
        RECT 57.530 178.350 57.760 178.690 ;
        RECT 66.170 178.630 66.400 178.690 ;
        RECT 67.190 178.630 67.420 178.690 ;
        RECT 66.170 178.350 67.420 178.630 ;
        RECT 75.830 178.350 76.060 178.690 ;
        RECT 57.530 178.090 76.060 178.350 ;
        RECT 57.530 177.700 57.760 178.090 ;
        RECT 66.170 177.790 67.420 178.090 ;
        RECT 66.170 177.700 66.400 177.790 ;
        RECT 67.190 177.730 67.420 177.790 ;
        RECT 75.830 177.730 76.060 178.090 ;
        RECT 57.530 177.440 66.400 177.700 ;
        RECT 67.630 177.680 75.610 177.700 ;
        RECT 67.625 177.450 75.625 177.680 ;
        RECT 67.630 177.440 75.610 177.450 ;
        RECT 76.360 177.080 79.600 179.310 ;
        RECT 85.380 179.160 85.680 179.860 ;
        RECT 86.080 179.360 86.380 179.660 ;
        RECT 85.900 179.160 86.130 179.210 ;
        RECT 85.380 178.260 86.130 179.160 ;
        RECT 85.900 178.210 86.130 178.260 ;
        RECT 86.340 179.160 86.570 179.210 ;
        RECT 87.480 179.160 87.780 179.860 ;
        RECT 88.180 179.360 88.480 179.660 ;
        RECT 88.000 179.160 88.230 179.210 ;
        RECT 86.340 178.260 86.980 179.160 ;
        RECT 87.480 178.260 88.230 179.160 ;
        RECT 86.340 178.210 86.570 178.260 ;
        RECT 27.070 176.720 79.600 177.080 ;
        RECT 80.130 177.360 81.280 177.630 ;
        RECT 86.080 177.360 86.380 178.060 ;
        RECT 80.130 176.960 86.380 177.360 ;
        RECT 86.080 176.260 86.380 176.960 ;
        RECT 86.780 177.360 86.980 178.260 ;
        RECT 88.000 178.210 88.230 178.260 ;
        RECT 88.440 179.160 88.670 179.210 ;
        RECT 88.440 178.260 89.080 179.160 ;
        RECT 88.440 178.210 88.670 178.260 ;
        RECT 88.180 177.360 88.480 178.060 ;
        RECT 86.780 176.960 88.480 177.360 ;
        RECT 34.985 175.870 44.985 176.100 ;
        RECT 34.550 175.760 34.780 175.820 ;
        RECT 45.190 175.760 45.420 175.820 ;
        RECT 34.480 174.920 34.840 175.760 ;
        RECT 45.120 174.920 45.480 175.760 ;
        RECT 34.550 174.860 34.780 174.920 ;
        RECT 45.190 174.860 45.420 174.920 ;
        RECT 34.995 174.810 44.975 174.840 ;
        RECT 34.985 174.580 44.985 174.810 ;
        RECT 24.460 173.740 25.190 174.510 ;
        RECT 51.010 174.430 51.740 176.170 ;
        RECT 61.905 175.870 71.905 176.100 ;
        RECT 85.900 176.060 86.130 176.065 ;
        RECT 61.470 175.760 61.700 175.820 ;
        RECT 72.110 175.760 72.340 175.820 ;
        RECT 61.400 174.920 61.760 175.760 ;
        RECT 72.040 174.920 72.400 175.760 ;
        RECT 61.470 174.860 61.700 174.920 ;
        RECT 72.110 174.860 72.340 174.920 ;
        RECT 61.915 174.810 71.895 174.840 ;
        RECT 61.905 174.580 71.905 174.810 ;
        RECT 51.010 174.140 54.290 174.430 ;
        RECT 53.950 173.740 54.290 174.140 ;
        RECT 85.380 174.160 86.130 176.060 ;
        RECT 24.460 173.480 51.370 173.740 ;
        RECT 53.950 173.480 78.290 173.740 ;
        RECT 24.460 172.480 25.190 173.480 ;
        RECT 38.480 172.830 39.200 172.870 ;
        RECT 40.560 172.830 41.260 172.840 ;
        RECT 29.195 172.600 39.200 172.830 ;
        RECT 40.555 172.600 50.550 172.830 ;
        RECT 38.480 172.550 39.200 172.600 ;
        RECT 40.560 172.570 41.650 172.600 ;
        RECT 28.740 172.490 29.020 172.550 ;
        RECT 28.390 172.300 29.020 172.490 ;
        RECT 28.390 170.090 28.580 172.300 ;
        RECT 28.740 172.240 29.020 172.300 ;
        RECT 39.380 172.240 39.650 172.550 ;
        RECT 40.100 172.240 40.380 172.550 ;
        RECT 50.740 172.490 51.010 172.550 ;
        RECT 51.180 172.490 51.370 173.480 ;
        RECT 65.400 172.830 66.120 172.870 ;
        RECT 67.480 172.830 68.180 172.840 ;
        RECT 56.115 172.600 66.120 172.830 ;
        RECT 67.475 172.600 77.470 172.830 ;
        RECT 65.400 172.550 66.120 172.600 ;
        RECT 67.480 172.570 68.570 172.600 ;
        RECT 55.660 172.490 55.940 172.550 ;
        RECT 50.740 172.300 51.370 172.490 ;
        RECT 50.740 172.240 51.010 172.300 ;
        RECT 29.220 172.190 29.940 172.230 ;
        RECT 40.550 172.190 41.650 172.200 ;
        RECT 49.810 172.190 50.530 172.240 ;
        RECT 29.195 171.960 39.190 172.190 ;
        RECT 40.550 171.960 50.550 172.190 ;
        RECT 29.220 171.910 29.940 171.960 ;
        RECT 40.550 171.940 41.650 171.960 ;
        RECT 49.810 171.900 50.530 171.960 ;
        RECT 38.480 171.630 39.200 171.670 ;
        RECT 40.560 171.630 41.280 171.680 ;
        RECT 29.195 171.400 39.200 171.630 ;
        RECT 40.555 171.400 50.550 171.630 ;
        RECT 38.480 171.350 39.200 171.400 ;
        RECT 28.720 171.040 29.040 171.350 ;
        RECT 39.340 171.020 39.680 171.370 ;
        RECT 40.070 171.020 40.410 171.370 ;
        RECT 40.560 171.350 41.280 171.400 ;
        RECT 50.710 171.020 51.040 171.380 ;
        RECT 30.420 170.990 31.140 171.020 ;
        RECT 48.610 170.990 49.330 171.000 ;
        RECT 29.195 170.760 39.190 170.990 ;
        RECT 40.555 170.760 50.550 170.990 ;
        RECT 30.420 170.710 31.140 170.760 ;
        RECT 48.610 170.740 49.330 170.760 ;
        RECT 38.480 170.430 39.200 170.470 ;
        RECT 40.560 170.430 41.280 170.480 ;
        RECT 29.195 170.200 39.200 170.430 ;
        RECT 40.555 170.200 50.550 170.430 ;
        RECT 38.480 170.150 39.200 170.200 ;
        RECT 40.560 170.170 41.610 170.200 ;
        RECT 28.740 170.090 29.020 170.150 ;
        RECT 28.390 169.900 29.020 170.090 ;
        RECT 28.390 167.790 28.580 169.900 ;
        RECT 28.740 169.840 29.020 169.900 ;
        RECT 39.380 169.840 39.650 170.150 ;
        RECT 40.100 169.840 40.380 170.150 ;
        RECT 50.740 170.090 51.010 170.150 ;
        RECT 51.180 170.090 51.370 172.300 ;
        RECT 50.740 169.900 51.370 170.090 ;
        RECT 55.310 172.300 55.940 172.490 ;
        RECT 55.310 170.090 55.500 172.300 ;
        RECT 55.660 172.240 55.940 172.300 ;
        RECT 66.300 172.240 66.570 172.550 ;
        RECT 67.020 172.240 67.300 172.550 ;
        RECT 77.660 172.490 77.930 172.550 ;
        RECT 78.100 172.490 78.290 173.480 ;
        RECT 85.380 173.370 85.680 174.160 ;
        RECT 85.900 174.065 86.130 174.160 ;
        RECT 86.340 176.060 86.570 176.065 ;
        RECT 86.780 176.060 86.980 176.960 ;
        RECT 88.180 176.260 88.480 176.960 ;
        RECT 88.880 177.360 89.080 178.260 ;
        RECT 88.880 176.960 89.280 177.360 ;
        RECT 88.000 176.060 88.230 176.065 ;
        RECT 86.340 174.160 86.980 176.060 ;
        RECT 87.480 174.160 88.230 176.060 ;
        RECT 86.340 174.065 86.570 174.160 ;
        RECT 86.080 173.560 86.380 173.860 ;
        RECT 87.480 173.370 87.780 174.160 ;
        RECT 88.000 174.065 88.230 174.160 ;
        RECT 88.440 176.060 88.670 176.065 ;
        RECT 88.880 176.060 89.080 176.960 ;
        RECT 88.440 174.160 89.080 176.060 ;
        RECT 88.440 174.065 88.670 174.160 ;
        RECT 88.180 173.560 88.480 173.860 ;
        RECT 85.180 172.570 104.140 173.370 ;
        RECT 77.660 172.300 78.290 172.490 ;
        RECT 77.660 172.240 77.930 172.300 ;
        RECT 56.140 172.190 56.860 172.230 ;
        RECT 67.470 172.190 68.570 172.200 ;
        RECT 76.730 172.190 77.450 172.240 ;
        RECT 56.115 171.960 66.110 172.190 ;
        RECT 67.470 171.960 77.470 172.190 ;
        RECT 56.140 171.910 56.860 171.960 ;
        RECT 67.470 171.940 68.570 171.960 ;
        RECT 76.730 171.900 77.450 171.960 ;
        RECT 65.400 171.630 66.120 171.670 ;
        RECT 67.480 171.630 68.200 171.680 ;
        RECT 56.115 171.400 66.120 171.630 ;
        RECT 67.475 171.400 77.470 171.630 ;
        RECT 65.400 171.350 66.120 171.400 ;
        RECT 55.640 171.040 55.960 171.350 ;
        RECT 66.260 171.020 66.600 171.370 ;
        RECT 66.990 171.020 67.330 171.370 ;
        RECT 67.480 171.350 68.200 171.400 ;
        RECT 77.630 171.020 77.960 171.380 ;
        RECT 57.340 170.990 58.060 171.020 ;
        RECT 75.530 170.990 76.250 171.000 ;
        RECT 56.115 170.760 66.110 170.990 ;
        RECT 67.475 170.760 77.470 170.990 ;
        RECT 57.340 170.710 58.060 170.760 ;
        RECT 75.530 170.740 76.250 170.760 ;
        RECT 65.400 170.430 66.120 170.470 ;
        RECT 67.480 170.430 68.200 170.480 ;
        RECT 56.115 170.200 66.120 170.430 ;
        RECT 67.475 170.200 77.470 170.430 ;
        RECT 65.400 170.150 66.120 170.200 ;
        RECT 67.480 170.170 68.530 170.200 ;
        RECT 55.660 170.090 55.940 170.150 ;
        RECT 55.310 169.900 55.940 170.090 ;
        RECT 50.740 169.840 51.010 169.900 ;
        RECT 29.220 169.790 29.940 169.830 ;
        RECT 40.550 169.790 41.610 169.800 ;
        RECT 49.810 169.790 50.530 169.840 ;
        RECT 29.195 169.560 39.190 169.790 ;
        RECT 40.550 169.560 50.550 169.790 ;
        RECT 29.220 169.510 29.940 169.560 ;
        RECT 40.550 169.540 41.610 169.560 ;
        RECT 49.810 169.500 50.530 169.560 ;
        RECT 38.480 169.230 39.200 169.270 ;
        RECT 40.560 169.230 41.280 169.280 ;
        RECT 29.195 169.000 39.200 169.230 ;
        RECT 40.555 169.000 50.550 169.230 ;
        RECT 38.480 168.950 39.200 169.000 ;
        RECT 28.720 168.640 29.040 168.950 ;
        RECT 39.340 168.620 39.680 168.970 ;
        RECT 40.070 168.620 40.410 168.970 ;
        RECT 40.560 168.950 41.280 169.000 ;
        RECT 50.710 168.620 51.040 168.980 ;
        RECT 30.420 168.590 31.140 168.620 ;
        RECT 48.610 168.590 49.330 168.600 ;
        RECT 29.195 168.360 39.190 168.590 ;
        RECT 40.555 168.360 50.550 168.590 ;
        RECT 30.420 168.310 31.140 168.360 ;
        RECT 48.610 168.340 49.330 168.360 ;
        RECT 52.980 167.790 53.620 168.800 ;
        RECT 55.310 167.790 55.500 169.900 ;
        RECT 55.660 169.840 55.940 169.900 ;
        RECT 66.300 169.840 66.570 170.150 ;
        RECT 67.020 169.840 67.300 170.150 ;
        RECT 77.660 170.090 77.930 170.150 ;
        RECT 78.100 170.090 78.290 172.300 ;
        RECT 77.660 169.900 78.290 170.090 ;
        RECT 85.380 171.780 85.680 172.570 ;
        RECT 86.080 172.080 86.380 172.380 ;
        RECT 85.900 171.780 86.130 171.875 ;
        RECT 77.660 169.840 77.930 169.900 ;
        RECT 85.380 169.880 86.130 171.780 ;
        RECT 85.900 169.875 86.130 169.880 ;
        RECT 86.340 171.780 86.570 171.875 ;
        RECT 87.480 171.780 87.780 172.570 ;
        RECT 88.180 172.080 88.480 172.380 ;
        RECT 88.000 171.780 88.230 171.875 ;
        RECT 86.340 169.880 86.980 171.780 ;
        RECT 87.480 169.880 88.230 171.780 ;
        RECT 86.340 169.875 86.570 169.880 ;
        RECT 56.140 169.790 56.860 169.830 ;
        RECT 67.470 169.790 68.530 169.800 ;
        RECT 76.730 169.790 77.450 169.840 ;
        RECT 56.115 169.560 66.110 169.790 ;
        RECT 67.470 169.560 77.470 169.790 ;
        RECT 56.140 169.510 56.860 169.560 ;
        RECT 67.470 169.540 68.530 169.560 ;
        RECT 76.730 169.500 77.450 169.560 ;
        RECT 65.400 169.230 66.120 169.270 ;
        RECT 67.480 169.230 68.200 169.280 ;
        RECT 56.115 169.000 66.120 169.230 ;
        RECT 67.475 169.000 77.470 169.230 ;
        RECT 65.400 168.950 66.120 169.000 ;
        RECT 55.640 168.640 55.960 168.950 ;
        RECT 66.260 168.620 66.600 168.970 ;
        RECT 66.990 168.620 67.330 168.970 ;
        RECT 67.480 168.950 68.200 169.000 ;
        RECT 86.080 168.980 86.380 169.680 ;
        RECT 77.630 168.620 77.960 168.980 ;
        RECT 57.340 168.590 58.060 168.620 ;
        RECT 75.530 168.590 76.250 168.600 ;
        RECT 56.115 168.360 66.110 168.590 ;
        RECT 67.475 168.360 77.470 168.590 ;
        RECT 83.780 168.580 86.380 168.980 ;
        RECT 57.340 168.310 58.060 168.360 ;
        RECT 75.530 168.340 76.250 168.360 ;
        RECT 83.780 168.100 84.740 168.580 ;
        RECT 86.080 167.880 86.380 168.580 ;
        RECT 86.780 168.980 86.980 169.880 ;
        RECT 88.000 169.875 88.230 169.880 ;
        RECT 88.440 171.780 88.670 171.875 ;
        RECT 88.440 169.880 89.080 171.780 ;
        RECT 88.440 169.875 88.670 169.880 ;
        RECT 88.180 168.980 88.480 169.680 ;
        RECT 86.780 168.580 88.480 168.980 ;
        RECT 20.500 167.530 51.040 167.790 ;
        RECT 52.980 167.530 77.960 167.790 ;
        RECT 85.900 167.680 86.130 167.730 ;
        RECT 20.500 165.760 22.660 167.530 ;
        RECT 30.410 167.130 50.530 167.390 ;
        RECT 29.210 166.730 49.330 166.990 ;
        RECT 52.980 166.420 53.620 167.530 ;
        RECT 57.330 167.130 77.450 167.390 ;
        RECT 56.130 166.730 76.250 166.990 ;
        RECT 85.380 166.780 86.130 167.680 ;
        RECT 85.380 166.080 85.680 166.780 ;
        RECT 85.900 166.730 86.130 166.780 ;
        RECT 86.340 167.680 86.570 167.730 ;
        RECT 86.780 167.680 86.980 168.580 ;
        RECT 88.180 167.880 88.480 168.580 ;
        RECT 88.880 168.980 89.080 169.880 ;
        RECT 88.880 168.580 89.280 168.980 ;
        RECT 88.000 167.680 88.230 167.730 ;
        RECT 86.340 166.780 86.980 167.680 ;
        RECT 87.480 166.780 88.230 167.680 ;
        RECT 86.340 166.730 86.570 166.780 ;
        RECT 86.080 166.280 86.380 166.580 ;
        RECT 87.480 166.080 87.780 166.780 ;
        RECT 88.000 166.730 88.230 166.780 ;
        RECT 88.440 167.680 88.670 167.730 ;
        RECT 88.880 167.680 89.080 168.580 ;
        RECT 88.440 166.780 89.080 167.680 ;
        RECT 88.440 166.730 88.670 166.780 ;
        RECT 88.180 166.280 88.480 166.580 ;
        RECT 27.730 165.850 32.110 165.870 ;
        RECT 33.980 165.850 38.960 165.870 ;
        RECT 40.950 165.850 45.930 165.870 ;
        RECT 27.730 165.610 32.510 165.850 ;
        RECT 33.970 165.620 38.970 165.850 ;
        RECT 40.940 165.620 45.940 165.850 ;
        RECT 33.980 165.610 38.960 165.620 ;
        RECT 40.950 165.610 45.930 165.620 ;
        RECT 47.270 165.610 52.020 165.870 ;
        RECT 27.730 165.220 27.960 165.610 ;
        RECT 32.280 165.510 32.510 165.610 ;
        RECT 47.270 165.590 47.630 165.610 ;
        RECT 47.270 165.570 47.470 165.590 ;
        RECT 33.580 165.510 33.810 165.570 ;
        RECT 39.130 165.510 39.360 165.570 ;
        RECT 40.550 165.510 40.780 165.570 ;
        RECT 46.100 165.510 46.330 165.570 ;
        RECT 47.240 165.510 47.470 165.570 ;
        RECT 32.280 165.220 33.810 165.510 ;
        RECT 39.060 165.220 39.420 165.510 ;
        RECT 27.730 164.960 39.420 165.220 ;
        RECT 12.770 144.800 14.930 157.770 ;
        RECT 20.500 145.180 22.660 164.630 ;
        RECT 27.730 164.610 27.960 164.960 ;
        RECT 32.280 164.670 33.810 164.960 ;
        RECT 39.060 164.670 39.420 164.960 ;
        RECT 40.490 165.220 40.850 165.510 ;
        RECT 46.100 165.220 47.470 165.510 ;
        RECT 51.790 165.220 52.020 165.610 ;
        RECT 40.490 164.960 52.020 165.220 ;
        RECT 40.490 164.670 40.850 164.960 ;
        RECT 46.100 164.670 47.470 164.960 ;
        RECT 32.280 164.610 32.510 164.670 ;
        RECT 33.580 164.610 33.810 164.670 ;
        RECT 39.130 164.610 39.360 164.670 ;
        RECT 40.550 164.610 40.780 164.670 ;
        RECT 46.100 164.610 46.330 164.670 ;
        RECT 47.240 164.610 47.470 164.670 ;
        RECT 51.790 164.610 52.020 164.960 ;
        RECT 54.650 165.850 59.030 165.870 ;
        RECT 60.900 165.850 65.880 165.870 ;
        RECT 67.870 165.850 72.850 165.870 ;
        RECT 54.650 165.610 59.430 165.850 ;
        RECT 60.890 165.620 65.890 165.850 ;
        RECT 67.860 165.620 72.860 165.850 ;
        RECT 60.900 165.610 65.880 165.620 ;
        RECT 67.870 165.610 72.850 165.620 ;
        RECT 74.190 165.610 78.940 165.870 ;
        RECT 54.650 165.220 54.880 165.610 ;
        RECT 59.200 165.510 59.430 165.610 ;
        RECT 74.190 165.590 74.550 165.610 ;
        RECT 74.190 165.570 74.390 165.590 ;
        RECT 60.500 165.510 60.730 165.570 ;
        RECT 66.050 165.510 66.280 165.570 ;
        RECT 67.470 165.510 67.700 165.570 ;
        RECT 73.020 165.510 73.250 165.570 ;
        RECT 74.160 165.510 74.390 165.570 ;
        RECT 59.200 165.220 60.730 165.510 ;
        RECT 65.980 165.220 66.340 165.510 ;
        RECT 54.650 164.960 66.340 165.220 ;
        RECT 54.650 164.610 54.880 164.960 ;
        RECT 59.200 164.670 60.730 164.960 ;
        RECT 65.980 164.670 66.340 164.960 ;
        RECT 67.410 165.220 67.770 165.510 ;
        RECT 73.020 165.220 74.390 165.510 ;
        RECT 78.710 165.220 78.940 165.610 ;
        RECT 85.180 165.450 104.140 166.080 ;
        RECT 67.410 164.960 78.940 165.220 ;
        RECT 67.410 164.670 67.770 164.960 ;
        RECT 73.020 164.670 74.390 164.960 ;
        RECT 59.200 164.610 59.430 164.670 ;
        RECT 60.500 164.610 60.730 164.670 ;
        RECT 66.050 164.610 66.280 164.670 ;
        RECT 67.470 164.610 67.700 164.670 ;
        RECT 73.020 164.610 73.250 164.670 ;
        RECT 74.160 164.610 74.390 164.670 ;
        RECT 78.710 164.610 78.940 164.960 ;
        RECT 28.120 164.330 32.120 164.560 ;
        RECT 33.970 164.330 38.970 164.560 ;
        RECT 40.940 164.330 45.940 164.560 ;
        RECT 47.630 164.330 51.630 164.560 ;
        RECT 55.040 164.330 59.040 164.560 ;
        RECT 60.890 164.330 65.890 164.560 ;
        RECT 67.860 164.330 72.860 164.560 ;
        RECT 74.550 164.330 78.550 164.560 ;
        RECT 28.430 163.960 31.800 164.330 ;
        RECT 34.720 163.960 38.090 164.330 ;
        RECT 41.830 163.960 45.200 164.330 ;
        RECT 55.350 163.960 58.720 164.330 ;
        RECT 61.640 163.960 65.010 164.330 ;
        RECT 68.750 163.960 72.120 164.330 ;
        RECT 89.080 163.970 104.140 165.450 ;
        RECT 85.180 163.960 104.140 163.970 ;
        RECT 27.070 163.790 104.140 163.960 ;
        RECT 27.070 161.560 32.990 163.790 ;
        RECT 33.980 163.420 38.960 163.440 ;
        RECT 40.950 163.420 45.930 163.440 ;
        RECT 33.970 163.190 38.970 163.420 ;
        RECT 40.940 163.190 45.940 163.420 ;
        RECT 33.980 163.180 38.960 163.190 ;
        RECT 40.950 163.180 45.930 163.190 ;
        RECT 33.580 162.800 33.810 163.140 ;
        RECT 39.130 163.080 39.360 163.140 ;
        RECT 40.550 163.080 40.780 163.140 ;
        RECT 39.060 162.800 39.420 163.080 ;
        RECT 33.580 162.540 39.420 162.800 ;
        RECT 33.580 162.180 33.810 162.540 ;
        RECT 39.060 162.240 39.420 162.540 ;
        RECT 40.490 162.800 40.850 163.080 ;
        RECT 46.100 162.800 46.330 163.140 ;
        RECT 40.490 162.540 46.330 162.800 ;
        RECT 40.490 162.240 40.850 162.540 ;
        RECT 39.130 162.180 39.360 162.240 ;
        RECT 40.550 162.180 40.780 162.240 ;
        RECT 46.100 162.180 46.330 162.540 ;
        RECT 33.970 161.900 38.970 162.130 ;
        RECT 40.940 161.900 45.940 162.130 ;
        RECT 34.030 161.560 38.910 161.900 ;
        RECT 41.000 161.560 45.880 161.900 ;
        RECT 46.760 161.560 59.910 163.790 ;
        RECT 60.900 163.420 65.880 163.440 ;
        RECT 67.870 163.420 72.850 163.440 ;
        RECT 60.890 163.190 65.890 163.420 ;
        RECT 67.860 163.190 72.860 163.420 ;
        RECT 60.900 163.180 65.880 163.190 ;
        RECT 67.870 163.180 72.850 163.190 ;
        RECT 60.500 162.800 60.730 163.140 ;
        RECT 66.050 163.080 66.280 163.140 ;
        RECT 67.470 163.080 67.700 163.140 ;
        RECT 65.980 162.800 66.340 163.080 ;
        RECT 60.500 162.540 66.340 162.800 ;
        RECT 60.500 162.180 60.730 162.540 ;
        RECT 65.980 162.240 66.340 162.540 ;
        RECT 67.410 162.800 67.770 163.080 ;
        RECT 73.020 162.800 73.250 163.140 ;
        RECT 67.410 162.540 73.250 162.800 ;
        RECT 67.410 162.240 67.770 162.540 ;
        RECT 66.050 162.180 66.280 162.240 ;
        RECT 67.470 162.180 67.700 162.240 ;
        RECT 73.020 162.180 73.250 162.540 ;
        RECT 60.890 161.900 65.890 162.130 ;
        RECT 67.860 161.900 72.860 162.130 ;
        RECT 60.950 161.560 65.830 161.900 ;
        RECT 67.920 161.560 72.800 161.900 ;
        RECT 73.680 161.560 104.140 163.790 ;
        RECT 27.070 160.800 104.140 161.560 ;
        RECT 27.070 159.460 59.910 160.800 ;
        RECT 60.950 160.460 65.830 160.800 ;
        RECT 67.920 160.460 72.800 160.800 ;
        RECT 60.890 160.230 65.890 160.460 ;
        RECT 67.860 160.230 72.860 160.460 ;
        RECT 44.810 159.120 49.690 159.460 ;
        RECT 44.750 158.890 49.750 159.120 ;
        RECT 44.360 158.780 44.590 158.840 ;
        RECT 49.910 158.780 50.140 158.840 ;
        RECT 43.700 157.860 44.590 158.780 ;
        RECT 44.750 157.810 49.750 157.830 ;
        RECT 49.890 157.810 50.190 158.780 ;
        RECT 53.990 158.570 59.910 159.460 ;
        RECT 60.500 159.820 60.730 160.180 ;
        RECT 66.050 160.120 66.280 160.180 ;
        RECT 67.470 160.120 67.700 160.180 ;
        RECT 65.980 159.820 66.340 160.120 ;
        RECT 60.500 159.560 66.340 159.820 ;
        RECT 60.500 159.220 60.730 159.560 ;
        RECT 65.980 159.280 66.340 159.560 ;
        RECT 67.410 159.820 67.770 160.120 ;
        RECT 73.020 159.820 73.250 160.180 ;
        RECT 67.410 159.560 73.250 159.820 ;
        RECT 67.410 159.280 67.770 159.560 ;
        RECT 66.050 159.220 66.280 159.280 ;
        RECT 67.470 159.220 67.700 159.280 ;
        RECT 73.020 159.220 73.250 159.560 ;
        RECT 60.900 159.170 65.880 159.180 ;
        RECT 67.870 159.170 72.850 159.180 ;
        RECT 60.890 158.940 65.890 159.170 ;
        RECT 67.860 158.940 72.860 159.170 ;
        RECT 60.900 158.920 65.880 158.940 ;
        RECT 67.870 158.920 72.850 158.940 ;
        RECT 73.680 158.570 104.140 160.800 ;
        RECT 53.990 158.400 104.140 158.570 ;
        RECT 55.350 158.030 58.720 158.400 ;
        RECT 61.640 158.030 65.010 158.400 ;
        RECT 68.750 158.030 72.120 158.400 ;
        RECT 44.750 157.600 50.190 157.810 ;
        RECT 55.040 157.800 59.040 158.030 ;
        RECT 60.890 157.800 65.890 158.030 ;
        RECT 67.860 157.800 72.860 158.030 ;
        RECT 74.550 157.800 78.550 158.030 ;
        RECT 38.810 152.190 40.970 156.140 ;
        RECT 47.810 154.730 50.190 157.600 ;
        RECT 54.650 157.400 54.880 157.750 ;
        RECT 59.200 157.690 59.430 157.750 ;
        RECT 60.500 157.690 60.730 157.750 ;
        RECT 66.050 157.690 66.280 157.750 ;
        RECT 67.470 157.690 67.700 157.750 ;
        RECT 73.020 157.690 73.250 157.750 ;
        RECT 74.160 157.690 74.390 157.750 ;
        RECT 59.200 157.400 60.730 157.690 ;
        RECT 65.980 157.400 66.340 157.690 ;
        RECT 54.650 157.140 66.340 157.400 ;
        RECT 54.650 156.750 54.880 157.140 ;
        RECT 59.200 156.850 60.730 157.140 ;
        RECT 65.980 156.850 66.340 157.140 ;
        RECT 67.410 157.400 67.770 157.690 ;
        RECT 73.020 157.400 74.390 157.690 ;
        RECT 78.710 157.400 78.940 157.750 ;
        RECT 67.410 157.140 78.940 157.400 ;
        RECT 67.410 156.850 67.770 157.140 ;
        RECT 73.020 156.850 74.390 157.140 ;
        RECT 59.200 156.750 59.430 156.850 ;
        RECT 60.500 156.790 60.730 156.850 ;
        RECT 66.050 156.790 66.280 156.850 ;
        RECT 67.470 156.790 67.700 156.850 ;
        RECT 73.020 156.790 73.250 156.850 ;
        RECT 74.160 156.790 74.390 156.850 ;
        RECT 74.190 156.770 74.390 156.790 ;
        RECT 74.190 156.750 74.550 156.770 ;
        RECT 78.710 156.750 78.940 157.140 ;
        RECT 54.650 156.510 59.430 156.750 ;
        RECT 60.900 156.740 65.880 156.750 ;
        RECT 67.870 156.740 72.850 156.750 ;
        RECT 60.890 156.510 65.890 156.740 ;
        RECT 67.860 156.510 72.860 156.740 ;
        RECT 54.650 156.490 59.030 156.510 ;
        RECT 60.900 156.490 65.880 156.510 ;
        RECT 67.870 156.490 72.850 156.510 ;
        RECT 74.190 156.490 78.940 156.750 ;
        RECT 52.770 154.830 53.500 155.920 ;
        RECT 56.130 155.370 76.250 155.630 ;
        RECT 57.330 154.970 77.450 155.230 ;
        RECT 52.770 154.570 77.960 154.830 ;
        RECT 24.420 147.750 25.730 150.080 ;
        RECT 38.810 147.110 40.970 151.060 ;
        RECT 47.810 149.650 49.970 153.600 ;
        RECT 52.770 153.480 53.500 154.570 ;
        RECT 55.310 152.460 55.500 154.570 ;
        RECT 57.340 154.000 58.060 154.050 ;
        RECT 75.530 154.000 76.250 154.020 ;
        RECT 56.115 153.770 66.110 154.000 ;
        RECT 67.475 153.770 77.470 154.000 ;
        RECT 57.340 153.740 58.060 153.770 ;
        RECT 75.530 153.760 76.250 153.770 ;
        RECT 55.640 153.410 55.960 153.720 ;
        RECT 65.400 153.360 66.120 153.410 ;
        RECT 66.260 153.390 66.600 153.740 ;
        RECT 66.990 153.390 67.330 153.740 ;
        RECT 67.480 153.360 68.200 153.410 ;
        RECT 77.630 153.380 77.960 153.740 ;
        RECT 56.115 153.130 66.120 153.360 ;
        RECT 67.475 153.130 77.470 153.360 ;
        RECT 65.400 153.090 66.120 153.130 ;
        RECT 67.480 153.080 68.200 153.130 ;
        RECT 56.140 152.800 56.860 152.850 ;
        RECT 67.470 152.800 68.530 152.820 ;
        RECT 76.730 152.800 77.450 152.860 ;
        RECT 56.115 152.570 66.110 152.800 ;
        RECT 67.470 152.570 77.470 152.800 ;
        RECT 56.140 152.530 56.860 152.570 ;
        RECT 67.470 152.560 68.530 152.570 ;
        RECT 76.730 152.520 77.450 152.570 ;
        RECT 55.660 152.460 55.940 152.520 ;
        RECT 55.310 152.270 55.940 152.460 ;
        RECT 55.310 150.060 55.500 152.270 ;
        RECT 55.660 152.210 55.940 152.270 ;
        RECT 66.300 152.210 66.570 152.520 ;
        RECT 67.020 152.210 67.300 152.520 ;
        RECT 77.660 152.460 77.930 152.520 ;
        RECT 77.660 152.270 78.290 152.460 ;
        RECT 77.660 152.210 77.930 152.270 ;
        RECT 65.400 152.160 66.120 152.210 ;
        RECT 67.480 152.160 68.530 152.190 ;
        RECT 56.115 151.930 66.120 152.160 ;
        RECT 67.475 151.930 77.470 152.160 ;
        RECT 65.400 151.890 66.120 151.930 ;
        RECT 67.480 151.880 68.200 151.930 ;
        RECT 57.340 151.600 58.060 151.650 ;
        RECT 75.530 151.600 76.250 151.620 ;
        RECT 56.115 151.370 66.110 151.600 ;
        RECT 67.475 151.370 77.470 151.600 ;
        RECT 57.340 151.340 58.060 151.370 ;
        RECT 75.530 151.360 76.250 151.370 ;
        RECT 55.640 151.010 55.960 151.320 ;
        RECT 65.400 150.960 66.120 151.010 ;
        RECT 66.260 150.990 66.600 151.340 ;
        RECT 66.990 150.990 67.330 151.340 ;
        RECT 67.480 150.960 68.200 151.010 ;
        RECT 77.630 150.980 77.960 151.340 ;
        RECT 56.115 150.730 66.120 150.960 ;
        RECT 67.475 150.730 77.470 150.960 ;
        RECT 65.400 150.690 66.120 150.730 ;
        RECT 67.480 150.680 68.200 150.730 ;
        RECT 56.140 150.400 56.860 150.450 ;
        RECT 67.470 150.400 68.570 150.420 ;
        RECT 76.730 150.400 77.450 150.460 ;
        RECT 56.115 150.170 66.110 150.400 ;
        RECT 67.470 150.170 77.470 150.400 ;
        RECT 56.140 150.130 56.860 150.170 ;
        RECT 67.470 150.160 68.570 150.170 ;
        RECT 76.730 150.120 77.450 150.170 ;
        RECT 55.660 150.060 55.940 150.120 ;
        RECT 55.310 149.870 55.940 150.060 ;
        RECT 55.660 149.810 55.940 149.870 ;
        RECT 66.300 149.810 66.570 150.120 ;
        RECT 67.020 149.810 67.300 150.120 ;
        RECT 77.660 150.060 77.930 150.120 ;
        RECT 78.100 150.060 78.290 152.270 ;
        RECT 77.660 149.870 78.290 150.060 ;
        RECT 77.660 149.810 77.930 149.870 ;
        RECT 65.400 149.760 66.120 149.810 ;
        RECT 67.480 149.760 68.570 149.790 ;
        RECT 56.115 149.530 66.120 149.760 ;
        RECT 67.475 149.530 77.470 149.760 ;
        RECT 65.400 149.490 66.120 149.530 ;
        RECT 67.480 149.520 68.180 149.530 ;
        RECT 50.980 148.880 53.060 149.090 ;
        RECT 78.100 148.880 78.290 149.870 ;
        RECT 50.980 148.620 78.290 148.880 ;
        RECT 34.170 144.880 36.190 146.650 ;
        RECT 47.810 145.310 49.970 148.520 ;
        RECT 50.980 148.410 53.060 148.620 ;
        RECT 61.905 147.550 71.905 147.780 ;
        RECT 61.915 147.520 71.895 147.550 ;
        RECT 61.470 147.440 61.700 147.500 ;
        RECT 72.110 147.440 72.340 147.500 ;
        RECT 61.400 146.600 61.760 147.440 ;
        RECT 72.040 146.600 72.400 147.440 ;
        RECT 61.470 146.540 61.700 146.600 ;
        RECT 72.110 146.540 72.340 146.600 ;
        RECT 61.905 146.260 71.905 146.490 ;
        RECT 47.810 145.230 50.660 145.310 ;
        RECT 39.445 145.030 50.660 145.230 ;
        RECT 39.445 145.000 49.445 145.030 ;
        RECT 38.530 144.880 39.300 144.970 ;
        RECT 11.930 142.070 23.490 144.800 ;
        RECT 34.170 144.020 39.300 144.880 ;
        RECT 49.620 144.380 50.660 145.030 ;
        RECT 53.990 145.280 104.120 145.640 ;
        RECT 49.620 144.050 49.970 144.380 ;
        RECT 39.005 143.990 39.235 144.020 ;
        RECT 49.655 143.990 49.885 144.050 ;
        RECT 39.445 143.920 49.445 143.940 ;
        RECT 39.430 143.700 49.460 143.920 ;
        RECT 53.990 143.700 57.230 145.280 ;
        RECT 27.070 143.050 57.230 143.700 ;
        RECT 57.530 144.660 66.400 144.920 ;
        RECT 67.630 144.910 75.610 144.920 ;
        RECT 67.625 144.680 75.625 144.910 ;
        RECT 67.630 144.660 75.610 144.680 ;
        RECT 57.530 144.270 57.760 144.660 ;
        RECT 66.170 144.570 66.400 144.660 ;
        RECT 67.190 144.570 67.420 144.630 ;
        RECT 66.170 144.270 67.420 144.570 ;
        RECT 75.830 144.270 76.060 144.630 ;
        RECT 57.530 144.010 76.060 144.270 ;
        RECT 57.530 143.670 57.760 144.010 ;
        RECT 66.170 143.730 67.420 144.010 ;
        RECT 66.170 143.670 66.400 143.730 ;
        RECT 67.190 143.670 67.420 143.730 ;
        RECT 75.830 143.670 76.060 144.010 ;
        RECT 57.965 143.390 65.965 143.620 ;
        RECT 67.625 143.390 75.625 143.620 ;
        RECT 58.025 143.050 65.905 143.390 ;
        RECT 67.685 143.050 75.565 143.390 ;
        RECT 76.350 143.050 104.120 145.280 ;
        RECT 27.070 142.040 104.120 143.050 ;
        RECT 27.070 142.030 79.600 142.040 ;
      LAYER met2 ;
        RECT 34.150 216.280 35.750 217.020 ;
        RECT 55.030 216.830 57.260 217.520 ;
        RECT 74.720 216.640 79.110 217.500 ;
        RECT 27.070 216.020 66.920 216.280 ;
        RECT 12.460 213.330 22.820 214.860 ;
        RECT 31.100 214.720 38.980 214.770 ;
        RECT 27.200 214.460 38.980 214.720 ;
        RECT 24.450 209.560 25.180 211.590 ;
        RECT 20.960 203.250 22.160 205.440 ;
        RECT 27.200 200.460 27.460 214.460 ;
        RECT 31.100 214.410 38.980 214.460 ;
        RECT 34.530 212.490 34.790 212.830 ;
        RECT 39.740 212.490 40.000 216.020 ;
        RECT 54.850 215.130 56.930 215.650 ;
        RECT 40.760 214.720 48.640 214.770 ;
        RECT 58.020 214.720 65.900 214.770 ;
        RECT 40.760 214.460 52.680 214.720 ;
        RECT 54.120 214.460 65.900 214.720 ;
        RECT 40.760 214.410 48.640 214.460 ;
        RECT 45.170 212.490 45.430 212.830 ;
        RECT 34.530 212.230 45.430 212.490 ;
        RECT 34.530 211.890 34.790 212.230 ;
        RECT 39.740 212.220 40.000 212.230 ;
        RECT 35.045 211.550 44.925 211.910 ;
        RECT 45.170 211.890 45.430 212.230 ;
        RECT 38.470 211.065 41.280 211.550 ;
        RECT 51.000 211.210 51.730 213.240 ;
        RECT 28.710 208.040 29.050 210.760 ;
        RECT 28.710 205.990 29.040 208.040 ;
        RECT 28.710 205.640 29.050 205.990 ;
        RECT 29.220 202.940 29.940 209.250 ;
        RECT 30.420 204.080 31.140 208.040 ;
        RECT 38.480 205.990 39.200 211.065 ;
        RECT 39.340 205.640 39.680 210.760 ;
        RECT 40.070 204.550 40.410 208.390 ;
        RECT 40.560 205.970 41.280 211.065 ;
        RECT 30.880 203.360 31.140 204.080 ;
        RECT 48.610 203.750 49.330 208.020 ;
        RECT 48.610 203.700 49.280 203.750 ;
        RECT 34.030 203.360 34.290 203.370 ;
        RECT 48.610 203.360 48.870 203.700 ;
        RECT 30.880 203.100 34.290 203.360 ;
        RECT 34.030 202.940 34.290 203.100 ;
        RECT 45.620 203.100 48.870 203.360 ;
        RECT 45.620 202.940 45.880 203.100 ;
        RECT 49.810 202.940 50.530 209.260 ;
        RECT 50.710 204.550 51.040 208.400 ;
        RECT 28.180 202.580 32.060 202.940 ;
        RECT 34.030 202.580 38.910 202.940 ;
        RECT 41.000 202.580 45.880 202.940 ;
        RECT 47.680 202.580 51.560 202.940 ;
        RECT 34.030 200.460 38.910 200.510 ;
        RECT 27.200 200.200 38.910 200.460 ;
        RECT 34.030 200.150 38.910 200.200 ;
        RECT 13.160 196.610 14.400 198.000 ;
        RECT 24.010 196.610 25.830 197.310 ;
        RECT 27.860 196.920 31.720 199.570 ;
        RECT 39.110 199.210 39.370 202.580 ;
        RECT 40.540 199.210 40.800 202.580 ;
        RECT 41.000 200.460 45.880 200.510 ;
        RECT 52.290 200.460 52.550 214.460 ;
        RECT 52.970 203.450 53.610 205.830 ;
        RECT 41.000 200.200 52.550 200.460 ;
        RECT 54.120 200.460 54.380 214.460 ;
        RECT 58.020 214.410 65.900 214.460 ;
        RECT 61.450 212.490 61.710 212.830 ;
        RECT 66.660 212.490 66.920 216.020 ;
        RECT 76.900 215.280 79.110 216.640 ;
        RECT 85.180 216.310 104.140 216.710 ;
        RECT 67.680 214.720 75.560 214.770 ;
        RECT 67.680 214.460 79.600 214.720 ;
        RECT 88.530 214.500 88.960 215.460 ;
        RECT 91.430 214.500 91.830 215.500 ;
        RECT 67.680 214.410 75.560 214.460 ;
        RECT 79.210 212.920 79.470 214.460 ;
        RECT 88.530 214.140 91.830 214.500 ;
        RECT 93.850 214.150 94.240 215.410 ;
        RECT 88.530 213.710 88.960 214.140 ;
        RECT 91.430 213.770 91.830 214.140 ;
        RECT 92.530 213.470 97.060 213.870 ;
        RECT 92.530 213.210 93.100 213.470 ;
        RECT 72.090 212.490 72.350 212.830 ;
        RECT 61.450 212.230 72.350 212.490 ;
        RECT 61.450 211.890 61.710 212.230 ;
        RECT 66.660 212.220 66.920 212.230 ;
        RECT 61.965 211.550 71.845 211.910 ;
        RECT 72.090 211.890 72.350 212.230 ;
        RECT 79.210 212.110 80.310 212.920 ;
        RECT 65.390 211.065 68.200 211.550 ;
        RECT 55.630 208.040 55.970 210.760 ;
        RECT 55.630 205.990 55.960 208.040 ;
        RECT 55.630 205.640 55.970 205.990 ;
        RECT 56.140 202.940 56.860 209.250 ;
        RECT 57.340 204.080 58.060 208.040 ;
        RECT 65.400 205.990 66.120 211.065 ;
        RECT 66.260 205.640 66.600 210.760 ;
        RECT 66.990 204.550 67.330 208.390 ;
        RECT 67.480 205.970 68.200 211.065 ;
        RECT 57.800 203.360 58.060 204.080 ;
        RECT 75.530 203.750 76.250 208.020 ;
        RECT 75.530 203.700 76.200 203.750 ;
        RECT 60.950 203.360 61.210 203.370 ;
        RECT 75.530 203.360 75.790 203.700 ;
        RECT 57.800 203.100 61.210 203.360 ;
        RECT 60.950 202.940 61.210 203.100 ;
        RECT 72.540 203.100 75.790 203.360 ;
        RECT 72.540 202.940 72.800 203.100 ;
        RECT 76.730 202.940 77.450 209.260 ;
        RECT 77.630 204.550 77.960 208.400 ;
        RECT 55.100 202.580 58.980 202.940 ;
        RECT 60.950 202.580 65.830 202.940 ;
        RECT 67.920 202.580 72.800 202.940 ;
        RECT 74.600 202.580 78.480 202.940 ;
        RECT 60.950 200.460 65.830 200.510 ;
        RECT 54.120 200.200 65.830 200.460 ;
        RECT 41.000 200.150 45.880 200.200 ;
        RECT 13.160 195.970 25.830 196.610 ;
        RECT 34.030 196.200 38.910 196.250 ;
        RECT 13.160 194.560 14.400 195.970 ;
        RECT 24.010 195.300 25.830 195.970 ;
        RECT 27.200 195.940 38.910 196.200 ;
        RECT 24.490 184.620 25.220 186.650 ;
        RECT 13.030 181.860 14.560 184.360 ;
        RECT 27.200 181.940 27.460 195.940 ;
        RECT 34.030 195.890 38.910 195.940 ;
        RECT 39.110 193.820 39.370 197.190 ;
        RECT 40.540 193.820 40.800 197.190 ;
        RECT 47.370 197.100 49.890 199.510 ;
        RECT 52.290 198.780 52.550 200.200 ;
        RECT 60.950 200.150 65.830 200.200 ;
        RECT 66.030 199.210 66.290 202.580 ;
        RECT 67.460 199.210 67.720 202.580 ;
        RECT 67.920 200.460 72.800 200.510 ;
        RECT 79.210 200.460 79.470 212.110 ;
        RECT 84.300 212.030 85.420 213.000 ;
        RECT 90.280 211.640 90.610 212.580 ;
        RECT 90.900 212.360 93.790 212.690 ;
        RECT 97.870 212.350 101.050 212.730 ;
        RECT 104.630 212.320 105.100 213.490 ;
        RECT 90.230 209.990 93.810 210.280 ;
        RECT 85.180 209.020 104.140 209.820 ;
        RECT 90.230 208.560 93.810 208.850 ;
        RECT 95.500 208.560 99.080 208.850 ;
        RECT 96.660 207.520 97.060 208.220 ;
        RECT 90.290 207.110 90.600 207.130 ;
        RECT 83.140 206.070 84.790 206.520 ;
        RECT 67.920 200.200 79.470 200.460 ;
        RECT 81.560 205.650 84.790 206.070 ;
        RECT 67.920 200.150 72.800 200.200 ;
        RECT 81.560 198.780 81.970 205.650 ;
        RECT 90.240 205.440 90.640 207.110 ;
        RECT 90.900 206.150 93.790 206.480 ;
        RECT 95.550 205.680 95.880 207.200 ;
        RECT 97.870 206.960 98.310 208.210 ;
        RECT 99.130 207.500 99.520 208.250 ;
        RECT 96.170 206.150 99.060 206.480 ;
        RECT 100.130 206.120 101.130 206.520 ;
        RECT 105.610 206.150 106.080 207.320 ;
        RECT 100.130 205.680 100.410 206.120 ;
        RECT 92.580 205.350 100.410 205.680 ;
        RECT 88.540 204.490 88.970 205.120 ;
        RECT 91.410 204.490 91.840 205.100 ;
        RECT 92.580 204.870 93.050 205.350 ;
        RECT 88.540 204.090 91.840 204.490 ;
        RECT 88.540 203.380 88.970 204.090 ;
        RECT 91.410 203.360 91.840 204.090 ;
        RECT 93.820 203.540 94.270 204.970 ;
        RECT 85.180 201.730 104.140 202.530 ;
        RECT 92.510 200.340 99.510 200.840 ;
        RECT 88.560 199.490 89.000 199.840 ;
        RECT 91.420 199.490 91.810 199.980 ;
        RECT 92.510 199.820 93.090 200.340 ;
        RECT 88.560 199.140 91.810 199.490 ;
        RECT 93.820 199.150 94.250 199.900 ;
        RECT 52.290 198.430 81.970 198.780 ;
        RECT 83.270 197.960 85.410 198.380 ;
        RECT 52.290 197.610 85.410 197.960 ;
        RECT 41.000 196.200 45.880 196.250 ;
        RECT 52.290 196.200 52.550 197.610 ;
        RECT 60.950 196.200 65.830 196.250 ;
        RECT 41.000 195.940 52.550 196.200 ;
        RECT 41.000 195.890 45.880 195.940 ;
        RECT 28.180 193.460 32.060 193.820 ;
        RECT 34.030 193.460 38.910 193.820 ;
        RECT 41.000 193.460 45.880 193.820 ;
        RECT 47.680 193.460 51.560 193.820 ;
        RECT 28.710 190.410 29.050 190.760 ;
        RECT 28.710 188.360 29.040 190.410 ;
        RECT 28.710 185.640 29.050 188.360 ;
        RECT 29.220 187.150 29.940 193.460 ;
        RECT 34.030 193.300 34.290 193.460 ;
        RECT 30.880 193.040 34.290 193.300 ;
        RECT 45.620 193.300 45.880 193.460 ;
        RECT 45.620 193.040 48.870 193.300 ;
        RECT 30.880 192.320 31.140 193.040 ;
        RECT 34.030 193.030 34.290 193.040 ;
        RECT 30.420 188.360 31.140 192.320 ;
        RECT 48.610 192.700 48.870 193.040 ;
        RECT 48.610 192.650 49.280 192.700 ;
        RECT 38.480 185.335 39.200 190.410 ;
        RECT 39.340 185.640 39.680 190.760 ;
        RECT 40.070 188.010 40.410 191.850 ;
        RECT 40.560 185.335 41.280 190.430 ;
        RECT 48.610 188.380 49.330 192.650 ;
        RECT 49.810 187.140 50.530 193.460 ;
        RECT 50.710 188.000 51.040 191.850 ;
        RECT 38.470 184.850 41.280 185.335 ;
        RECT 34.530 184.170 34.790 184.510 ;
        RECT 35.045 184.490 44.925 184.850 ;
        RECT 39.740 184.170 40.000 184.180 ;
        RECT 45.170 184.170 45.430 184.510 ;
        RECT 34.530 183.910 45.430 184.170 ;
        RECT 34.530 183.570 34.790 183.910 ;
        RECT 31.100 181.940 38.980 181.990 ;
        RECT 27.200 181.680 38.980 181.940 ;
        RECT 31.100 181.630 38.980 181.680 ;
        RECT 39.740 180.380 40.000 183.910 ;
        RECT 45.170 183.570 45.430 183.910 ;
        RECT 51.080 183.140 51.810 185.170 ;
        RECT 40.760 181.940 48.640 181.990 ;
        RECT 52.290 181.940 52.550 195.940 ;
        RECT 54.120 195.940 65.830 196.200 ;
        RECT 53.000 190.440 53.640 192.820 ;
        RECT 54.120 181.940 54.380 195.940 ;
        RECT 60.950 195.890 65.830 195.940 ;
        RECT 66.030 193.820 66.290 197.190 ;
        RECT 67.460 193.820 67.720 197.190 ;
        RECT 90.280 196.720 90.610 198.820 ;
        RECT 90.900 197.780 93.790 198.110 ;
        RECT 98.720 197.280 99.400 198.230 ;
        RECT 107.100 197.760 107.570 198.930 ;
        RECT 98.720 196.720 99.050 197.280 ;
        RECT 90.280 196.380 99.050 196.720 ;
        RECT 67.920 196.200 72.800 196.250 ;
        RECT 67.920 195.940 79.470 196.200 ;
        RECT 67.920 195.890 72.800 195.940 ;
        RECT 55.100 193.460 58.980 193.820 ;
        RECT 60.950 193.460 65.830 193.820 ;
        RECT 67.920 193.460 72.800 193.820 ;
        RECT 74.600 193.460 78.480 193.820 ;
        RECT 55.630 190.410 55.970 190.760 ;
        RECT 55.630 188.360 55.960 190.410 ;
        RECT 55.630 185.640 55.970 188.360 ;
        RECT 56.140 187.150 56.860 193.460 ;
        RECT 60.950 193.300 61.210 193.460 ;
        RECT 57.800 193.040 61.210 193.300 ;
        RECT 72.540 193.300 72.800 193.460 ;
        RECT 72.540 193.040 75.790 193.300 ;
        RECT 57.800 192.320 58.060 193.040 ;
        RECT 60.950 193.030 61.210 193.040 ;
        RECT 57.340 188.360 58.060 192.320 ;
        RECT 75.530 192.700 75.790 193.040 ;
        RECT 75.530 192.650 76.200 192.700 ;
        RECT 65.400 185.335 66.120 190.410 ;
        RECT 66.260 185.640 66.600 190.760 ;
        RECT 66.990 188.010 67.330 191.850 ;
        RECT 67.480 185.335 68.200 190.430 ;
        RECT 75.530 188.380 76.250 192.650 ;
        RECT 76.730 187.140 77.450 193.460 ;
        RECT 79.210 192.100 79.470 195.940 ;
        RECT 90.230 195.410 93.810 195.700 ;
        RECT 85.180 194.440 104.140 195.240 ;
        RECT 90.000 193.430 90.890 194.100 ;
        RECT 77.630 188.000 77.960 191.850 ;
        RECT 79.210 191.410 79.980 192.100 ;
        RECT 65.390 184.850 68.200 185.335 ;
        RECT 61.450 184.170 61.710 184.510 ;
        RECT 61.965 184.490 71.845 184.850 ;
        RECT 66.660 184.170 66.920 184.180 ;
        RECT 72.090 184.170 72.350 184.510 ;
        RECT 61.450 183.910 72.350 184.170 ;
        RECT 61.450 183.570 61.710 183.910 ;
        RECT 58.020 181.940 65.900 181.990 ;
        RECT 40.760 181.680 52.680 181.940 ;
        RECT 54.120 181.680 65.900 181.940 ;
        RECT 40.760 181.630 48.640 181.680 ;
        RECT 58.020 181.630 65.900 181.680 ;
        RECT 54.730 180.720 56.750 181.350 ;
        RECT 66.660 180.380 66.920 183.910 ;
        RECT 72.090 183.570 72.350 183.910 ;
        RECT 67.680 181.940 75.560 181.990 ;
        RECT 79.210 181.940 79.470 191.410 ;
        RECT 82.410 191.240 83.520 192.260 ;
        RECT 85.180 187.150 104.140 187.950 ;
        RECT 88.560 185.670 88.970 186.210 ;
        RECT 93.070 185.670 93.460 186.270 ;
        RECT 88.560 185.260 93.460 185.670 ;
        RECT 88.560 184.640 88.970 185.260 ;
        RECT 81.570 182.920 83.430 183.870 ;
        RECT 180.310 183.560 183.110 183.840 ;
        RECT 180.310 183.280 183.390 183.560 ;
        RECT 180.310 183.000 183.670 183.280 ;
        RECT 67.680 181.680 79.600 181.940 ;
        RECT 67.680 181.630 75.560 181.680 ;
        RECT 27.070 179.010 66.920 180.380 ;
        RECT 27.070 179.000 40.000 179.010 ;
        RECT 53.990 179.000 66.920 179.010 ;
        RECT 31.100 177.700 38.980 177.750 ;
        RECT 27.200 177.440 38.980 177.700 ;
        RECT 24.460 172.480 25.190 174.510 ;
        RECT 13.270 166.240 14.550 168.580 ;
        RECT 27.200 163.440 27.460 177.440 ;
        RECT 31.100 177.390 38.980 177.440 ;
        RECT 34.530 175.470 34.790 175.810 ;
        RECT 39.740 175.470 40.000 179.000 ;
        RECT 54.670 177.990 56.820 178.610 ;
        RECT 40.760 177.700 48.640 177.750 ;
        RECT 58.020 177.700 65.900 177.750 ;
        RECT 40.760 177.440 52.680 177.700 ;
        RECT 54.120 177.440 65.900 177.700 ;
        RECT 40.760 177.390 48.640 177.440 ;
        RECT 45.170 175.470 45.430 175.810 ;
        RECT 34.530 175.210 45.430 175.470 ;
        RECT 34.530 174.870 34.790 175.210 ;
        RECT 39.740 175.200 40.000 175.210 ;
        RECT 35.045 174.530 44.925 174.890 ;
        RECT 45.170 174.870 45.430 175.210 ;
        RECT 38.470 174.045 41.280 174.530 ;
        RECT 51.010 174.140 51.740 176.170 ;
        RECT 28.710 171.020 29.050 173.740 ;
        RECT 28.710 168.970 29.040 171.020 ;
        RECT 28.710 168.620 29.050 168.970 ;
        RECT 29.220 165.920 29.940 172.230 ;
        RECT 30.420 167.060 31.140 171.020 ;
        RECT 38.480 168.970 39.200 174.045 ;
        RECT 39.340 168.620 39.680 173.740 ;
        RECT 40.070 167.530 40.410 171.370 ;
        RECT 40.560 168.950 41.280 174.045 ;
        RECT 30.880 166.340 31.140 167.060 ;
        RECT 48.610 166.730 49.330 171.000 ;
        RECT 48.610 166.680 49.280 166.730 ;
        RECT 34.030 166.340 34.290 166.350 ;
        RECT 48.610 166.340 48.870 166.680 ;
        RECT 30.880 166.080 34.290 166.340 ;
        RECT 34.030 165.920 34.290 166.080 ;
        RECT 45.620 166.080 48.870 166.340 ;
        RECT 45.620 165.920 45.880 166.080 ;
        RECT 49.810 165.920 50.530 172.240 ;
        RECT 50.710 167.530 51.040 171.380 ;
        RECT 28.180 165.560 32.060 165.920 ;
        RECT 34.030 165.560 38.910 165.920 ;
        RECT 41.000 165.560 45.880 165.920 ;
        RECT 47.680 165.560 51.560 165.920 ;
        RECT 34.030 163.440 38.910 163.490 ;
        RECT 27.200 163.180 38.910 163.440 ;
        RECT 34.030 163.130 38.910 163.180 ;
        RECT 27.570 159.750 31.430 162.400 ;
        RECT 39.110 162.190 39.370 165.560 ;
        RECT 40.540 162.190 40.800 165.560 ;
        RECT 41.000 163.440 45.880 163.490 ;
        RECT 52.290 163.440 52.550 177.440 ;
        RECT 52.980 166.420 53.620 168.800 ;
        RECT 41.000 163.180 52.550 163.440 ;
        RECT 54.120 163.440 54.380 177.440 ;
        RECT 58.020 177.390 65.900 177.440 ;
        RECT 61.450 175.470 61.710 175.810 ;
        RECT 66.660 175.470 66.920 179.000 ;
        RECT 76.830 178.540 79.150 180.990 ;
        RECT 67.680 177.700 75.560 177.750 ;
        RECT 67.680 177.440 81.320 177.700 ;
        RECT 67.680 177.390 75.560 177.440 ;
        RECT 79.210 177.140 81.320 177.440 ;
        RECT 72.090 175.470 72.350 175.810 ;
        RECT 61.450 175.210 72.350 175.470 ;
        RECT 61.450 174.870 61.710 175.210 ;
        RECT 66.660 175.200 66.920 175.210 ;
        RECT 61.965 174.530 71.845 174.890 ;
        RECT 72.090 174.870 72.350 175.210 ;
        RECT 65.390 174.045 68.200 174.530 ;
        RECT 55.630 171.020 55.970 173.740 ;
        RECT 55.630 168.970 55.960 171.020 ;
        RECT 55.630 168.620 55.970 168.970 ;
        RECT 56.140 165.920 56.860 172.230 ;
        RECT 57.340 167.060 58.060 171.020 ;
        RECT 65.400 168.970 66.120 174.045 ;
        RECT 66.260 168.620 66.600 173.740 ;
        RECT 66.990 167.530 67.330 171.370 ;
        RECT 67.480 168.950 68.200 174.045 ;
        RECT 57.800 166.340 58.060 167.060 ;
        RECT 75.530 166.730 76.250 171.000 ;
        RECT 75.530 166.680 76.200 166.730 ;
        RECT 60.950 166.340 61.210 166.350 ;
        RECT 75.530 166.340 75.790 166.680 ;
        RECT 57.800 166.080 61.210 166.340 ;
        RECT 60.950 165.920 61.210 166.080 ;
        RECT 72.540 166.080 75.790 166.340 ;
        RECT 72.540 165.920 72.800 166.080 ;
        RECT 76.730 165.920 77.450 172.240 ;
        RECT 77.630 167.530 77.960 171.380 ;
        RECT 55.100 165.560 58.980 165.920 ;
        RECT 60.950 165.560 65.830 165.920 ;
        RECT 67.920 165.560 72.800 165.920 ;
        RECT 74.600 165.560 78.480 165.920 ;
        RECT 60.950 163.440 65.830 163.490 ;
        RECT 54.120 163.180 65.830 163.440 ;
        RECT 41.000 163.130 45.880 163.180 ;
        RECT 47.410 160.280 49.680 162.610 ;
        RECT 52.290 161.400 52.550 163.180 ;
        RECT 60.950 163.130 65.830 163.180 ;
        RECT 66.030 162.190 66.290 165.560 ;
        RECT 67.460 162.190 67.720 165.560 ;
        RECT 67.920 163.440 72.800 163.490 ;
        RECT 79.210 163.440 79.470 177.140 ;
        RECT 67.920 163.180 79.470 163.440 ;
        RECT 67.920 163.130 72.800 163.180 ;
        RECT 82.270 161.400 82.700 182.920 ;
        RECT 180.310 182.720 181.150 183.000 ;
        RECT 182.550 182.720 183.670 183.000 ;
        RECT 184.790 182.720 185.630 183.840 ;
        RECT 189.270 183.280 190.670 183.840 ;
        RECT 188.990 183.000 190.670 183.280 ;
        RECT 188.990 182.720 189.550 183.000 ;
        RECT 180.030 182.440 181.150 182.720 ;
        RECT 147.550 181.600 149.230 181.880 ;
        RECT 146.710 181.320 149.230 181.600 ;
        RECT 180.030 181.320 180.870 182.440 ;
        RECT 182.830 182.160 183.670 182.720 ;
        RECT 184.510 182.440 185.630 182.720 ;
        RECT 146.150 181.040 149.230 181.320 ;
        RECT 145.870 180.760 149.230 181.040 ;
        RECT 85.180 179.860 104.140 180.660 ;
        RECT 145.590 179.920 148.950 180.760 ;
        RECT 179.750 180.200 180.590 181.320 ;
        RECT 182.550 180.760 183.390 182.160 ;
        RECT 184.510 181.320 185.350 182.440 ;
        RECT 188.710 181.880 189.550 182.720 ;
        RECT 182.270 180.480 183.110 180.760 ;
        RECT 181.990 180.200 183.110 180.480 ;
        RECT 154.830 179.920 156.790 180.200 ;
        RECT 179.750 179.920 182.830 180.200 ;
        RECT 184.230 179.920 185.070 181.320 ;
        RECT 188.430 181.040 189.270 181.880 ;
        RECT 188.150 180.480 188.990 181.040 ;
        RECT 189.830 180.480 190.670 183.000 ;
        RECT 192.630 182.720 193.470 183.840 ;
        RECT 195.430 183.560 196.550 183.840 ;
        RECT 197.110 183.560 199.910 183.840 ;
        RECT 195.430 183.280 196.270 183.560 ;
        RECT 195.150 183.000 195.990 183.280 ;
        RECT 192.350 182.440 193.470 182.720 ;
        RECT 194.870 182.720 195.990 183.000 ;
        RECT 197.110 183.000 199.630 183.560 ;
        RECT 197.110 182.720 197.950 183.000 ;
        RECT 202.710 182.720 204.390 183.840 ;
        RECT 206.350 183.280 208.030 183.840 ;
        RECT 209.990 183.560 211.950 183.840 ;
        RECT 213.630 183.700 216.710 183.840 ;
        RECT 213.630 183.560 216.570 183.700 ;
        RECT 216.990 183.560 220.070 183.840 ;
        RECT 209.710 183.280 212.230 183.560 ;
        RECT 194.870 182.440 195.710 182.720 ;
        RECT 196.830 182.440 197.950 182.720 ;
        RECT 192.350 181.320 193.190 182.440 ;
        RECT 194.590 181.880 195.430 182.440 ;
        RECT 194.310 181.600 195.150 181.880 ;
        RECT 194.030 181.320 195.150 181.600 ;
        RECT 196.830 181.320 197.670 182.440 ;
        RECT 202.430 181.320 203.270 182.720 ;
        RECT 203.830 182.440 204.390 182.720 ;
        RECT 206.070 182.720 208.030 183.280 ;
        RECT 209.150 183.000 212.230 183.280 ;
        RECT 213.350 183.000 216.430 183.560 ;
        RECT 216.710 183.000 219.790 183.560 ;
        RECT 209.150 182.720 210.270 183.000 ;
        RECT 206.070 182.440 206.630 182.720 ;
        RECT 188.150 180.200 188.710 180.480 ;
        RECT 189.830 180.200 190.390 180.480 ;
        RECT 145.310 177.680 148.950 179.920 ;
        RECT 154.270 179.640 155.110 179.920 ;
        RECT 153.990 179.360 154.550 179.640 ;
        RECT 156.510 179.360 156.790 179.920 ;
        RECT 153.430 179.080 154.270 179.360 ;
        RECT 156.230 179.080 156.790 179.360 ;
        RECT 179.470 179.360 182.550 179.920 ;
        RECT 153.150 178.800 153.710 179.080 ;
        RECT 155.950 178.800 156.510 179.080 ;
        RECT 179.470 178.800 180.310 179.360 ;
        RECT 181.710 179.080 182.830 179.360 ;
        RECT 152.590 178.520 153.430 178.800 ;
        RECT 155.670 178.520 156.230 178.800 ;
        RECT 179.190 178.520 180.310 178.800 ;
        RECT 181.990 178.800 183.110 179.080 ;
        RECT 183.950 178.800 184.790 179.920 ;
        RECT 187.870 179.640 188.710 180.200 ;
        RECT 187.590 178.800 188.430 179.640 ;
        RECT 152.310 178.240 152.870 178.520 ;
        RECT 155.390 178.240 155.950 178.520 ;
        RECT 152.030 177.960 152.590 178.240 ;
        RECT 154.830 177.960 155.670 178.240 ;
        RECT 151.470 177.680 152.310 177.960 ;
        RECT 154.550 177.680 155.390 177.960 ;
        RECT 145.030 177.400 148.950 177.680 ;
        RECT 151.190 177.400 151.750 177.680 ;
        RECT 154.270 177.400 154.830 177.680 ;
        RECT 179.190 177.400 180.030 178.520 ;
        RECT 181.990 177.680 182.830 178.800 ;
        RECT 183.670 178.520 184.790 178.800 ;
        RECT 187.310 178.520 188.150 178.800 ;
        RECT 189.550 178.520 190.390 180.200 ;
        RECT 192.070 180.200 192.910 181.320 ;
        RECT 194.030 181.040 194.870 181.320 ;
        RECT 193.750 180.480 194.590 181.040 ;
        RECT 193.470 180.200 194.310 180.480 ;
        RECT 196.550 180.200 197.390 181.320 ;
        RECT 192.070 179.920 194.030 180.200 ;
        RECT 196.550 179.920 198.790 180.200 ;
        RECT 202.150 179.920 202.990 181.320 ;
        RECT 203.550 181.040 204.390 182.440 ;
        RECT 205.790 181.880 206.630 182.440 ;
        RECT 205.790 181.600 206.350 181.880 ;
        RECT 206.910 181.600 207.750 182.720 ;
        RECT 208.870 182.440 209.990 182.720 ;
        RECT 208.870 181.600 209.710 182.440 ;
        RECT 205.510 181.040 206.350 181.600 ;
        RECT 191.790 179.360 194.030 179.920 ;
        RECT 191.790 178.800 192.630 179.360 ;
        RECT 83.520 176.960 84.800 177.360 ;
        RECT 145.030 176.280 148.670 177.400 ;
        RECT 150.910 177.120 151.470 177.400 ;
        RECT 153.990 177.120 154.550 177.400 ;
        RECT 150.630 176.840 151.190 177.120 ;
        RECT 153.710 176.840 154.270 177.120 ;
        RECT 150.350 176.560 150.910 176.840 ;
        RECT 153.430 176.560 153.990 176.840 ;
        RECT 149.790 176.280 150.630 176.560 ;
        RECT 153.150 176.280 153.710 176.560 ;
        RECT 145.030 176.000 148.110 176.280 ;
        RECT 149.510 176.000 150.070 176.280 ;
        RECT 152.870 176.000 153.430 176.280 ;
        RECT 88.540 175.260 88.990 175.860 ;
        RECT 145.030 175.720 147.550 176.000 ;
        RECT 149.230 175.720 149.790 176.000 ;
        RECT 152.310 175.720 153.150 176.000 ;
        RECT 144.750 175.440 146.990 175.720 ;
        RECT 148.950 175.440 149.510 175.720 ;
        RECT 152.030 175.440 152.870 175.720 ;
        RECT 88.540 174.840 92.650 175.260 ;
        RECT 144.750 174.880 146.430 175.440 ;
        RECT 148.670 175.160 149.230 175.440 ;
        RECT 151.750 175.160 152.590 175.440 ;
        RECT 159.310 175.160 163.230 176.840 ;
        RECT 178.910 176.280 179.750 177.400 ;
        RECT 181.710 176.560 182.550 177.680 ;
        RECT 183.670 177.400 184.510 178.520 ;
        RECT 187.310 177.960 190.390 178.520 ;
        RECT 187.030 177.680 190.390 177.960 ;
        RECT 181.150 176.280 182.550 176.560 ;
        RECT 183.390 176.280 184.230 177.400 ;
        RECT 187.030 177.120 187.870 177.680 ;
        RECT 186.750 176.560 187.590 177.120 ;
        RECT 186.470 176.280 187.590 176.560 ;
        RECT 189.550 176.280 190.390 177.680 ;
        RECT 191.510 178.520 192.630 178.800 ;
        RECT 193.190 178.800 194.030 179.360 ;
        RECT 196.270 179.360 198.790 179.920 ;
        RECT 196.270 178.800 197.110 179.360 ;
        RECT 201.870 178.800 202.710 179.920 ;
        RECT 203.550 179.360 204.110 181.040 ;
        RECT 205.510 180.760 206.070 181.040 ;
        RECT 205.230 180.200 206.070 180.760 ;
        RECT 206.630 180.200 207.470 181.600 ;
        RECT 208.590 181.320 209.710 181.600 ;
        RECT 211.390 182.160 212.510 183.000 ;
        RECT 214.470 182.160 215.310 183.000 ;
        RECT 217.830 182.160 218.670 183.000 ;
        RECT 208.590 180.200 209.430 181.320 ;
        RECT 211.390 181.040 212.230 182.160 ;
        RECT 214.190 181.040 215.030 182.160 ;
        RECT 217.550 181.040 218.390 182.160 ;
        RECT 205.230 179.920 205.790 180.200 ;
        RECT 191.510 177.400 192.350 178.520 ;
        RECT 193.190 178.240 194.310 178.800 ;
        RECT 193.470 177.400 194.310 178.240 ;
        RECT 195.990 178.520 197.110 178.800 ;
        RECT 201.590 178.520 202.710 178.800 ;
        RECT 195.990 177.400 196.830 178.520 ;
        RECT 201.590 177.400 202.430 178.520 ;
        RECT 203.270 177.960 204.110 179.360 ;
        RECT 204.950 179.360 205.790 179.920 ;
        RECT 204.950 179.080 205.510 179.360 ;
        RECT 206.350 179.080 207.190 180.200 ;
        RECT 204.670 178.520 205.510 179.080 ;
        RECT 206.070 178.800 207.190 179.080 ;
        RECT 208.310 178.800 209.150 180.200 ;
        RECT 211.110 179.640 211.950 181.040 ;
        RECT 213.910 180.760 215.030 181.040 ;
        RECT 217.270 180.760 218.390 181.040 ;
        RECT 213.910 179.640 214.750 180.760 ;
        RECT 217.270 179.640 218.110 180.760 ;
        RECT 204.670 178.240 205.230 178.520 ;
        RECT 178.910 176.000 182.270 176.280 ;
        RECT 183.390 176.000 185.910 176.280 ;
        RECT 178.630 175.720 181.990 176.000 ;
        RECT 178.630 175.440 181.430 175.720 ;
        RECT 183.110 175.440 185.630 176.000 ;
        RECT 186.470 175.720 187.310 176.280 ;
        RECT 189.270 175.720 190.390 176.280 ;
        RECT 191.230 176.000 192.070 177.400 ;
        RECT 193.470 176.840 194.590 177.400 ;
        RECT 193.750 176.000 194.590 176.840 ;
        RECT 195.710 176.280 196.550 177.400 ;
        RECT 195.710 176.000 198.230 176.280 ;
        RECT 201.310 176.000 202.150 177.400 ;
        RECT 203.270 176.280 203.830 177.960 ;
        RECT 204.390 177.680 205.230 178.240 ;
        RECT 206.070 177.680 206.910 178.800 ;
        RECT 208.030 177.680 208.870 178.800 ;
        RECT 210.830 178.520 211.670 179.640 ;
        RECT 204.390 177.400 204.950 177.680 ;
        RECT 204.110 176.840 204.950 177.400 ;
        RECT 204.110 176.280 204.670 176.840 ;
        RECT 205.790 176.280 206.630 177.680 ;
        RECT 207.750 177.400 208.870 177.680 ;
        RECT 210.550 178.240 211.670 178.520 ;
        RECT 213.630 179.360 214.750 179.640 ;
        RECT 216.990 179.360 218.110 179.640 ;
        RECT 213.630 178.240 214.470 179.360 ;
        RECT 216.990 178.240 217.830 179.360 ;
        RECT 207.750 176.560 208.590 177.400 ;
        RECT 210.550 177.120 211.390 178.240 ;
        RECT 210.270 176.840 211.390 177.120 ;
        RECT 213.350 176.840 214.190 178.240 ;
        RECT 216.710 176.840 217.550 178.240 ;
        RECT 210.270 176.560 211.110 176.840 ;
        RECT 207.750 176.280 208.870 176.560 ;
        RECT 209.990 176.280 211.110 176.560 ;
        RECT 202.990 176.000 204.670 176.280 ;
        RECT 186.190 175.440 187.030 175.720 ;
        RECT 189.270 175.440 190.110 175.720 ;
        RECT 190.950 175.440 191.790 176.000 ;
        RECT 193.750 175.440 194.870 176.000 ;
        RECT 195.430 175.440 198.230 176.000 ;
        RECT 201.030 175.440 201.870 176.000 ;
        RECT 202.990 175.440 204.390 176.000 ;
        RECT 205.510 175.440 206.350 176.280 ;
        RECT 207.750 176.000 210.830 176.280 ;
        RECT 208.030 175.720 210.550 176.000 ;
        RECT 213.070 175.720 213.910 176.840 ;
        RECT 216.430 175.720 217.270 176.840 ;
        RECT 208.310 175.440 210.270 175.720 ;
        RECT 212.790 175.440 213.910 175.720 ;
        RECT 216.150 175.440 217.270 175.720 ;
        RECT 148.390 174.880 148.950 175.160 ;
        RECT 151.470 174.880 152.310 175.160 ;
        RECT 159.310 174.880 163.510 175.160 ;
        RECT 88.540 174.290 88.990 174.840 ;
        RECT 144.750 174.600 146.150 174.880 ;
        RECT 148.110 174.600 148.670 174.880 ;
        RECT 151.190 174.600 152.030 174.880 ;
        RECT 159.310 174.600 165.750 174.880 ;
        RECT 144.470 174.320 146.150 174.600 ;
        RECT 147.830 174.320 148.390 174.600 ;
        RECT 150.910 174.320 151.470 174.600 ;
        RECT 159.310 174.320 166.310 174.600 ;
        RECT 144.470 174.040 145.870 174.320 ;
        RECT 147.550 174.040 148.110 174.320 ;
        RECT 150.630 174.040 151.470 174.320 ;
        RECT 159.030 174.040 167.150 174.320 ;
        RECT 144.190 173.480 145.870 174.040 ;
        RECT 147.270 173.760 147.830 174.040 ;
        RECT 150.350 173.760 150.910 174.040 ;
        RECT 151.330 173.900 151.750 174.040 ;
        RECT 146.990 173.480 147.550 173.760 ;
        RECT 150.070 173.480 150.630 173.760 ;
        RECT 151.470 173.480 151.750 173.900 ;
        RECT 159.030 173.760 167.710 174.040 ;
        RECT 159.030 173.480 168.270 173.760 ;
        RECT 85.180 172.570 104.140 173.370 ;
        RECT 144.190 172.640 145.590 173.480 ;
        RECT 146.710 173.200 147.270 173.480 ;
        RECT 149.510 173.200 150.350 173.480 ;
        RECT 151.610 173.340 152.030 173.480 ;
        RECT 146.430 172.920 146.990 173.200 ;
        RECT 149.230 172.920 150.070 173.200 ;
        RECT 151.750 172.920 152.030 173.340 ;
        RECT 158.750 173.200 168.830 173.480 ;
        RECT 158.750 172.920 169.390 173.200 ;
        RECT 178.070 172.920 217.830 173.760 ;
        RECT 146.150 172.640 146.710 172.920 ;
        RECT 148.950 172.640 149.790 172.920 ;
        RECT 151.750 172.640 152.310 172.920 ;
        RECT 143.910 172.360 146.430 172.640 ;
        RECT 148.670 172.360 149.510 172.640 ;
        RECT 88.530 170.480 88.960 171.590 ;
        RECT 143.910 171.520 146.150 172.360 ;
        RECT 148.110 172.080 149.230 172.360 ;
        RECT 152.030 172.080 152.310 172.640 ;
        RECT 158.470 172.640 169.950 172.920 ;
        RECT 158.470 172.360 170.790 172.640 ;
        RECT 177.790 172.360 217.550 172.920 ;
        RECT 158.190 172.080 171.350 172.360 ;
        RECT 147.830 171.800 148.950 172.080 ;
        RECT 152.170 171.940 152.590 172.080 ;
        RECT 146.990 171.520 148.950 171.800 ;
        RECT 152.310 171.800 152.590 171.940 ;
        RECT 158.190 171.800 171.910 172.080 ;
        RECT 177.790 171.800 217.270 172.360 ;
        RECT 152.310 171.520 152.870 171.800 ;
        RECT 143.910 171.240 147.830 171.520 ;
        RECT 143.910 170.960 147.270 171.240 ;
        RECT 148.390 170.960 148.950 171.520 ;
        RECT 152.590 171.240 152.870 171.520 ;
        RECT 157.910 171.520 164.630 171.800 ;
        RECT 165.750 171.520 172.470 171.800 ;
        RECT 177.790 171.520 216.990 171.800 ;
        RECT 157.910 171.240 164.350 171.520 ;
        RECT 166.590 171.240 172.470 171.520 ;
        RECT 152.590 170.960 153.150 171.240 ;
        RECT 88.530 170.040 94.220 170.480 ;
        RECT 144.190 170.400 147.550 170.960 ;
        RECT 148.390 170.400 149.230 170.960 ;
        RECT 152.870 170.680 153.150 170.960 ;
        RECT 157.630 170.960 164.350 171.240 ;
        RECT 167.710 170.960 172.470 171.240 ;
        RECT 157.630 170.680 164.070 170.960 ;
        RECT 168.830 170.680 172.470 170.960 ;
        RECT 153.010 170.540 153.430 170.680 ;
        RECT 143.910 170.120 147.270 170.400 ;
        RECT 148.670 170.120 149.510 170.400 ;
        RECT 153.150 170.120 153.430 170.540 ;
        RECT 157.350 170.120 164.070 170.680 ;
        RECT 169.670 170.400 172.190 170.680 ;
        RECT 143.630 169.560 147.270 170.120 ;
        RECT 148.950 169.840 149.790 170.120 ;
        RECT 153.290 169.980 153.710 170.120 ;
        RECT 143.350 169.280 143.910 169.560 ;
        RECT 144.190 169.280 147.270 169.560 ;
        RECT 149.230 169.560 150.070 169.840 ;
        RECT 153.430 169.560 153.710 169.980 ;
        RECT 157.070 169.560 163.790 170.120 ;
        RECT 149.230 169.280 150.630 169.560 ;
        RECT 153.570 169.420 153.990 169.560 ;
        RECT 153.710 169.280 153.990 169.420 ;
        RECT 143.070 169.000 143.630 169.280 ;
        RECT 144.190 169.000 146.990 169.280 ;
        RECT 149.790 169.000 151.190 169.280 ;
        RECT 153.710 169.000 154.270 169.280 ;
        RECT 156.790 169.000 164.070 169.560 ;
        RECT 52.290 161.040 82.700 161.400 ;
        RECT 83.780 168.100 84.740 168.970 ;
        RECT 142.790 168.440 143.350 169.000 ;
        RECT 144.470 168.720 146.990 169.000 ;
        RECT 150.070 168.720 152.030 169.000 ;
        RECT 153.990 168.720 154.270 169.000 ;
        RECT 144.470 168.440 146.710 168.720 ;
        RECT 150.630 168.440 153.150 168.720 ;
        RECT 154.130 168.580 154.550 168.720 ;
        RECT 154.270 168.440 154.550 168.580 ;
        RECT 156.510 168.440 164.350 169.000 ;
        RECT 173.030 168.720 179.750 169.000 ;
        RECT 169.670 168.440 186.750 168.720 ;
        RECT 142.510 168.160 143.070 168.440 ;
        RECT 144.470 168.160 146.430 168.440 ;
        RECT 151.470 168.160 154.830 168.440 ;
        RECT 60.950 159.180 65.830 159.230 ;
        RECT 54.120 158.920 65.830 159.180 ;
        RECT 20.650 155.230 22.260 155.820 ;
        RECT 52.770 155.230 53.500 155.920 ;
        RECT 20.650 154.520 53.500 155.230 ;
        RECT 20.650 153.880 22.260 154.520 ;
        RECT 52.770 153.480 53.500 154.520 ;
        RECT 24.420 149.090 25.730 150.080 ;
        RECT 24.420 148.410 53.060 149.090 ;
        RECT 24.420 147.750 25.730 148.410 ;
        RECT 34.170 144.850 36.190 146.650 ;
        RECT 11.930 142.070 23.490 144.800 ;
        RECT 49.620 144.380 50.660 145.310 ;
        RECT 54.120 144.920 54.380 158.920 ;
        RECT 60.950 158.870 65.830 158.920 ;
        RECT 66.030 156.800 66.290 160.170 ;
        RECT 67.460 156.800 67.720 160.170 ;
        RECT 67.920 159.180 72.800 159.230 ;
        RECT 83.780 159.180 84.220 168.100 ;
        RECT 142.230 167.600 142.790 168.160 ;
        RECT 144.470 167.880 146.150 168.160 ;
        RECT 152.310 167.880 155.110 168.160 ;
        RECT 156.230 167.880 164.350 168.440 ;
        RECT 168.830 168.160 189.550 168.440 ;
        RECT 168.270 167.880 170.510 168.160 ;
        RECT 185.630 167.880 190.950 168.160 ;
        RECT 144.750 167.600 145.870 167.880 ;
        RECT 153.430 167.600 164.350 167.880 ;
        RECT 167.710 167.600 169.390 167.880 ;
        RECT 188.990 167.600 191.510 167.880 ;
        RECT 141.950 167.040 142.510 167.600 ;
        RECT 154.270 167.320 164.350 167.600 ;
        RECT 167.430 167.320 168.550 167.600 ;
        RECT 190.670 167.320 191.790 167.600 ;
        RECT 143.910 167.040 144.190 167.320 ;
        RECT 155.110 167.040 164.070 167.320 ;
        RECT 167.150 167.040 168.270 167.320 ;
        RECT 191.230 167.040 192.070 167.320 ;
        RECT 141.670 166.480 142.230 167.040 ;
        RECT 143.630 166.760 144.190 167.040 ;
        RECT 155.950 166.760 164.070 167.040 ;
        RECT 166.870 166.760 167.710 167.040 ;
        RECT 191.510 166.760 192.350 167.040 ;
        RECT 143.630 166.480 143.910 166.760 ;
        RECT 149.790 166.480 150.070 166.760 ;
        RECT 156.790 166.480 164.070 166.760 ;
        RECT 166.590 166.480 167.430 166.760 ;
        RECT 191.790 166.480 192.630 166.760 ;
        RECT 85.180 165.680 104.140 166.080 ;
        RECT 141.390 165.920 141.950 166.480 ;
        RECT 143.350 166.340 143.770 166.480 ;
        RECT 143.350 166.200 143.630 166.340 ;
        RECT 149.230 166.200 150.070 166.480 ;
        RECT 157.630 166.200 163.790 166.480 ;
        RECT 166.310 166.200 167.150 166.480 ;
        RECT 143.070 165.920 143.630 166.200 ;
        RECT 148.950 165.920 149.790 166.200 ;
        RECT 158.190 165.920 163.790 166.200 ;
        RECT 166.030 165.920 166.870 166.200 ;
        RECT 187.310 165.920 190.670 166.200 ;
        RECT 192.070 165.920 192.910 166.480 ;
        RECT 100.520 164.950 103.170 165.680 ;
        RECT 141.110 165.360 141.670 165.920 ;
        RECT 143.070 165.640 143.350 165.920 ;
        RECT 148.390 165.640 149.510 165.920 ;
        RECT 159.030 165.640 163.790 165.920 ;
        RECT 140.830 165.080 141.670 165.360 ;
        RECT 142.790 165.360 143.350 165.640 ;
        RECT 148.110 165.360 148.950 165.640 ;
        RECT 159.870 165.360 163.790 165.640 ;
        RECT 165.750 165.360 166.590 165.920 ;
        RECT 176.670 165.640 180.590 165.920 ;
        RECT 185.630 165.640 191.510 165.920 ;
        RECT 192.350 165.640 193.190 165.920 ;
        RECT 174.710 165.360 177.510 165.640 ;
        RECT 184.230 165.360 187.310 165.640 ;
        RECT 190.110 165.360 191.790 165.640 ;
        RECT 192.630 165.360 193.470 165.640 ;
        RECT 142.790 165.080 143.070 165.360 ;
        RECT 147.830 165.080 148.670 165.360 ;
        RECT 160.710 165.080 163.510 165.360 ;
        RECT 165.470 165.080 166.310 165.360 ;
        RECT 173.310 165.080 175.830 165.360 ;
        RECT 183.110 165.080 185.630 165.360 ;
        RECT 190.950 165.080 192.070 165.360 ;
        RECT 192.910 165.080 193.750 165.360 ;
        RECT 140.830 164.520 141.390 165.080 ;
        RECT 142.510 164.800 143.070 165.080 ;
        RECT 147.270 164.800 148.390 165.080 ;
        RECT 161.550 164.800 164.350 165.080 ;
        RECT 165.470 164.800 166.030 165.080 ;
        RECT 171.910 164.800 174.430 165.080 ;
        RECT 181.990 164.800 184.230 165.080 ;
        RECT 191.230 164.800 192.070 165.080 ;
        RECT 193.190 164.800 194.030 165.080 ;
        RECT 142.510 164.520 142.790 164.800 ;
        RECT 146.990 164.520 147.830 164.800 ;
        RECT 162.670 164.520 166.030 164.800 ;
        RECT 170.790 164.520 173.310 164.800 ;
        RECT 181.150 164.520 182.830 164.800 ;
        RECT 191.510 164.520 192.070 164.800 ;
        RECT 193.470 164.520 194.030 164.800 ;
        RECT 140.550 163.680 141.110 164.520 ;
        RECT 142.230 164.240 142.790 164.520 ;
        RECT 146.710 164.240 147.550 164.520 ;
        RECT 163.510 164.240 166.870 164.520 ;
        RECT 169.670 164.240 172.190 164.520 ;
        RECT 180.310 164.240 181.710 164.520 ;
        RECT 142.230 163.960 142.510 164.240 ;
        RECT 146.430 163.960 147.270 164.240 ;
        RECT 164.630 163.960 171.070 164.240 ;
        RECT 179.470 163.960 180.870 164.240 ;
        RECT 140.270 163.400 141.110 163.680 ;
        RECT 141.950 163.400 142.510 163.960 ;
        RECT 146.150 163.680 146.990 163.960 ;
        RECT 166.030 163.680 169.950 163.960 ;
        RECT 178.630 163.680 180.030 163.960 ;
        RECT 191.510 163.680 192.350 164.520 ;
        RECT 193.470 164.240 194.310 164.520 ;
        RECT 193.750 163.960 194.590 164.240 ;
        RECT 194.030 163.680 194.870 163.960 ;
        RECT 145.870 163.400 146.710 163.680 ;
        RECT 165.750 163.400 167.990 163.680 ;
        RECT 168.550 163.400 169.670 163.680 ;
        RECT 178.070 163.400 179.190 163.680 ;
        RECT 191.790 163.400 192.630 163.680 ;
        RECT 194.310 163.400 194.870 163.680 ;
        RECT 140.270 162.560 140.830 163.400 ;
        RECT 141.950 163.120 142.230 163.400 ;
        RECT 145.590 163.120 146.430 163.400 ;
        RECT 164.910 163.120 167.150 163.400 ;
        RECT 168.830 163.120 169.950 163.400 ;
        RECT 177.230 163.120 178.350 163.400 ;
        RECT 191.790 163.120 192.910 163.400 ;
        RECT 194.310 163.120 195.150 163.400 ;
        RECT 141.670 162.560 142.230 163.120 ;
        RECT 145.310 162.840 146.150 163.120 ;
        RECT 163.790 162.840 166.310 163.120 ;
        RECT 169.110 162.840 170.230 163.120 ;
        RECT 176.670 162.840 177.510 163.120 ;
        RECT 192.070 162.840 192.910 163.120 ;
        RECT 194.590 162.840 195.430 163.120 ;
        RECT 145.030 162.560 145.870 162.840 ;
        RECT 162.950 162.560 165.190 162.840 ;
        RECT 169.390 162.560 170.510 162.840 ;
        RECT 176.670 162.560 176.950 162.840 ;
        RECT 192.070 162.560 193.190 162.840 ;
        RECT 194.870 162.560 195.710 162.840 ;
        RECT 139.990 162.280 140.830 162.560 ;
        RECT 139.990 160.880 140.550 162.280 ;
        RECT 141.390 161.720 141.950 162.560 ;
        RECT 145.030 162.280 145.590 162.560 ;
        RECT 162.110 162.280 164.350 162.560 ;
        RECT 169.950 162.280 170.790 162.560 ;
        RECT 192.350 162.280 193.470 162.560 ;
        RECT 195.150 162.280 195.710 162.560 ;
        RECT 144.750 162.000 145.310 162.280 ;
        RECT 161.270 162.000 163.510 162.280 ;
        RECT 170.230 162.000 171.350 162.280 ;
        RECT 192.630 162.000 193.750 162.280 ;
        RECT 195.150 162.000 195.990 162.280 ;
        RECT 144.470 161.720 145.310 162.000 ;
        RECT 160.430 161.720 162.670 162.000 ;
        RECT 170.510 161.720 171.630 162.000 ;
        RECT 192.910 161.720 194.310 162.000 ;
        RECT 195.430 161.720 196.270 162.000 ;
        RECT 141.390 161.440 141.670 161.720 ;
        RECT 67.920 158.920 84.220 159.180 ;
        RECT 139.710 159.760 140.550 160.880 ;
        RECT 141.110 160.320 141.670 161.440 ;
        RECT 144.190 161.440 145.030 161.720 ;
        RECT 159.590 161.440 161.550 161.720 ;
        RECT 170.790 161.440 171.910 161.720 ;
        RECT 193.190 161.440 194.590 161.720 ;
        RECT 195.150 161.440 196.270 161.720 ;
        RECT 144.190 161.160 144.750 161.440 ;
        RECT 158.470 161.160 160.710 161.440 ;
        RECT 171.070 161.160 172.470 161.440 ;
        RECT 193.470 161.160 196.550 161.440 ;
        RECT 143.910 160.880 144.750 161.160 ;
        RECT 157.630 160.880 159.870 161.160 ;
        RECT 171.630 160.880 173.030 161.160 ;
        RECT 193.750 160.880 195.710 161.160 ;
        RECT 195.990 160.880 196.830 161.160 ;
        RECT 143.910 160.600 144.470 160.880 ;
        RECT 156.790 160.600 159.030 160.880 ;
        RECT 171.910 160.600 173.590 160.880 ;
        RECT 193.750 160.600 195.150 160.880 ;
        RECT 196.270 160.600 197.110 160.880 ;
        RECT 143.630 160.320 144.190 160.600 ;
        RECT 155.950 160.320 158.190 160.600 ;
        RECT 172.470 160.320 174.150 160.600 ;
        RECT 193.190 160.320 194.590 160.600 ;
        RECT 196.550 160.320 197.110 160.600 ;
        RECT 67.920 158.870 72.800 158.920 ;
        RECT 55.100 156.440 58.980 156.800 ;
        RECT 60.950 156.440 65.830 156.800 ;
        RECT 67.920 156.440 72.800 156.800 ;
        RECT 74.600 156.440 78.480 156.800 ;
        RECT 55.630 153.390 55.970 153.740 ;
        RECT 55.630 151.340 55.960 153.390 ;
        RECT 55.630 148.620 55.970 151.340 ;
        RECT 56.140 150.130 56.860 156.440 ;
        RECT 60.950 156.280 61.210 156.440 ;
        RECT 57.800 156.020 61.210 156.280 ;
        RECT 72.540 156.280 72.800 156.440 ;
        RECT 72.540 156.020 75.790 156.280 ;
        RECT 57.800 155.300 58.060 156.020 ;
        RECT 60.950 156.010 61.210 156.020 ;
        RECT 57.340 151.340 58.060 155.300 ;
        RECT 75.530 155.680 75.790 156.020 ;
        RECT 75.530 155.630 76.200 155.680 ;
        RECT 65.400 148.315 66.120 153.390 ;
        RECT 66.260 148.620 66.600 153.740 ;
        RECT 66.990 150.990 67.330 154.830 ;
        RECT 67.480 148.315 68.200 153.410 ;
        RECT 75.530 151.360 76.250 155.630 ;
        RECT 76.730 150.120 77.450 156.440 ;
        RECT 77.630 150.980 77.960 154.830 ;
        RECT 65.390 147.830 68.200 148.315 ;
        RECT 61.450 147.150 61.710 147.490 ;
        RECT 61.965 147.470 71.845 147.830 ;
        RECT 66.660 147.150 66.920 147.160 ;
        RECT 72.090 147.150 72.350 147.490 ;
        RECT 61.450 146.890 72.350 147.150 ;
        RECT 61.450 146.550 61.710 146.890 ;
        RECT 58.020 144.920 65.900 144.970 ;
        RECT 54.120 144.660 65.900 144.920 ;
        RECT 58.020 144.610 65.900 144.660 ;
        RECT 50.230 143.360 50.660 144.380 ;
        RECT 54.710 143.700 56.860 144.320 ;
        RECT 66.660 143.360 66.920 146.890 ;
        RECT 72.090 146.550 72.350 146.890 ;
        RECT 67.680 144.920 75.560 144.970 ;
        RECT 79.210 144.920 79.470 158.920 ;
        RECT 139.710 158.080 140.270 159.760 ;
        RECT 139.710 157.240 140.550 158.080 ;
        RECT 140.830 157.240 141.390 160.320 ;
        RECT 143.350 160.040 144.190 160.320 ;
        RECT 155.110 160.040 157.350 160.320 ;
        RECT 167.710 160.040 168.270 160.320 ;
        RECT 173.030 160.040 174.430 160.320 ;
        RECT 192.910 160.040 194.310 160.320 ;
        RECT 196.830 160.040 197.390 160.320 ;
        RECT 143.350 159.760 143.910 160.040 ;
        RECT 154.270 159.760 156.510 160.040 ;
        RECT 167.150 159.760 167.990 160.040 ;
        RECT 173.590 159.760 174.430 160.040 ;
        RECT 192.630 159.760 193.750 160.040 ;
        RECT 196.830 159.760 197.670 160.040 ;
        RECT 143.070 159.480 143.910 159.760 ;
        RECT 153.430 159.480 155.670 159.760 ;
        RECT 166.310 159.480 167.430 159.760 ;
        RECT 173.870 159.480 174.430 159.760 ;
        RECT 192.070 159.480 193.470 159.760 ;
        RECT 197.110 159.480 197.670 159.760 ;
        RECT 143.070 158.920 143.630 159.480 ;
        RECT 152.590 159.200 154.830 159.480 ;
        RECT 165.750 159.200 166.870 159.480 ;
        RECT 151.750 158.920 153.710 159.200 ;
        RECT 142.790 158.360 143.350 158.920 ;
        RECT 150.910 158.640 152.870 158.920 ;
        RECT 150.070 158.360 152.030 158.640 ;
        RECT 142.510 158.080 143.350 158.360 ;
        RECT 149.230 158.080 151.190 158.360 ;
        RECT 142.510 157.520 143.070 158.080 ;
        RECT 148.390 157.800 150.350 158.080 ;
        RECT 147.550 157.520 149.510 157.800 ;
        RECT 154.550 157.520 154.830 159.200 ;
        RECT 164.910 158.920 166.310 159.200 ;
        RECT 172.190 158.920 172.750 159.200 ;
        RECT 173.870 158.920 174.710 159.480 ;
        RECT 191.790 159.200 192.910 159.480 ;
        RECT 197.390 159.200 197.950 159.480 ;
        RECT 191.510 158.920 192.630 159.200 ;
        RECT 164.350 158.640 165.470 158.920 ;
        RECT 171.630 158.640 172.470 158.920 ;
        RECT 163.510 158.360 164.910 158.640 ;
        RECT 171.070 158.360 172.190 158.640 ;
        RECT 162.950 158.080 164.350 158.360 ;
        RECT 170.510 158.080 171.910 158.360 ;
        RECT 174.150 158.080 174.710 158.920 ;
        RECT 191.230 158.640 192.350 158.920 ;
        RECT 197.670 158.640 198.230 159.200 ;
        RECT 190.950 158.360 192.070 158.640 ;
        RECT 197.950 158.360 198.510 158.640 ;
        RECT 162.110 157.800 163.790 158.080 ;
        RECT 169.950 157.800 171.630 158.080 ;
        RECT 161.550 157.520 163.230 157.800 ;
        RECT 169.670 157.520 171.350 157.800 ;
        RECT 139.710 156.680 141.390 157.240 ;
        RECT 142.230 157.240 143.070 157.520 ;
        RECT 146.710 157.240 148.670 157.520 ;
        RECT 153.990 157.380 154.690 157.520 ;
        RECT 153.990 157.240 154.550 157.380 ;
        RECT 160.710 157.240 162.670 157.520 ;
        RECT 169.110 157.240 171.070 157.520 ;
        RECT 139.990 156.400 141.670 156.680 ;
        RECT 142.230 156.400 142.790 157.240 ;
        RECT 145.870 156.960 147.830 157.240 ;
        RECT 153.710 156.960 154.270 157.240 ;
        RECT 160.150 156.960 162.110 157.240 ;
        RECT 168.550 156.960 170.790 157.240 ;
        RECT 145.030 156.680 146.990 156.960 ;
        RECT 153.150 156.820 153.850 156.960 ;
        RECT 153.150 156.680 153.710 156.820 ;
        RECT 159.310 156.680 161.550 156.960 ;
        RECT 167.990 156.680 170.510 156.960 ;
        RECT 174.150 156.680 174.990 158.080 ;
        RECT 190.950 157.800 191.790 158.360 ;
        RECT 198.230 158.080 198.790 158.360 ;
        RECT 191.230 157.240 192.070 157.800 ;
        RECT 198.510 157.520 199.070 158.080 ;
        RECT 198.790 157.240 199.350 157.520 ;
        RECT 191.510 156.960 192.350 157.240 ;
        RECT 199.070 156.960 199.630 157.240 ;
        RECT 191.790 156.680 192.630 156.960 ;
        RECT 144.190 156.400 146.150 156.680 ;
        RECT 146.710 156.400 147.270 156.680 ;
        RECT 152.590 156.540 153.290 156.680 ;
        RECT 152.590 156.400 153.150 156.540 ;
        RECT 158.750 156.400 160.710 156.680 ;
        RECT 167.430 156.400 170.230 156.680 ;
        RECT 140.550 156.120 142.790 156.400 ;
        RECT 143.350 156.120 145.310 156.400 ;
        RECT 146.990 156.120 147.270 156.400 ;
        RECT 152.030 156.260 152.730 156.400 ;
        RECT 152.030 156.120 152.590 156.260 ;
        RECT 158.190 156.120 160.150 156.400 ;
        RECT 166.870 156.120 168.270 156.400 ;
        RECT 168.830 156.120 169.950 156.400 ;
        RECT 174.150 156.120 174.710 156.680 ;
        RECT 192.070 156.400 192.910 156.680 ;
        RECT 192.350 156.120 193.190 156.400 ;
        RECT 206.070 156.120 206.630 156.400 ;
        RECT 140.830 155.840 144.750 156.120 ;
        RECT 147.130 155.980 147.550 156.120 ;
        RECT 147.270 155.840 147.550 155.980 ;
        RECT 151.470 155.980 152.170 156.120 ;
        RECT 151.470 155.840 152.030 155.980 ;
        RECT 157.350 155.840 159.590 156.120 ;
        RECT 166.310 155.840 167.710 156.120 ;
        RECT 168.830 155.840 169.670 156.120 ;
        RECT 173.870 155.840 174.990 156.120 ;
        RECT 192.630 155.840 193.470 156.120 ;
        RECT 205.790 155.840 206.910 156.120 ;
        RECT 141.390 155.560 143.910 155.840 ;
        RECT 147.270 155.560 147.830 155.840 ;
        RECT 150.630 155.700 151.610 155.840 ;
        RECT 150.630 155.560 151.470 155.700 ;
        RECT 156.790 155.560 159.030 155.840 ;
        RECT 165.750 155.560 167.150 155.840 ;
        RECT 168.830 155.560 169.390 155.840 ;
        RECT 173.590 155.560 175.270 155.840 ;
        RECT 192.910 155.560 193.750 155.840 ;
        RECT 205.510 155.560 207.190 155.840 ;
        RECT 141.670 155.280 143.350 155.560 ;
        RECT 147.550 155.280 148.110 155.560 ;
        RECT 150.070 155.280 150.910 155.560 ;
        RECT 155.950 155.280 158.470 155.560 ;
        RECT 165.470 155.280 166.590 155.560 ;
        RECT 168.550 155.280 169.110 155.560 ;
        RECT 173.590 155.280 174.430 155.560 ;
        RECT 174.990 155.280 175.830 155.560 ;
        RECT 193.190 155.280 194.030 155.560 ;
        RECT 204.950 155.280 206.630 155.560 ;
        RECT 141.950 155.000 143.910 155.280 ;
        RECT 147.970 155.140 150.210 155.280 ;
        RECT 148.110 155.000 150.070 155.140 ;
        RECT 155.390 155.000 157.910 155.280 ;
        RECT 164.910 155.000 166.030 155.280 ;
        RECT 168.270 155.000 168.830 155.280 ;
        RECT 173.590 155.000 174.150 155.280 ;
        RECT 175.550 155.000 176.110 155.280 ;
        RECT 192.630 155.000 194.310 155.280 ;
        RECT 204.670 155.000 206.350 155.280 ;
        RECT 206.910 155.000 207.190 155.560 ;
        RECT 142.510 154.720 144.190 155.000 ;
        RECT 154.550 154.720 157.350 155.000 ;
        RECT 164.350 154.720 165.470 155.000 ;
        RECT 167.990 154.720 168.550 155.000 ;
        RECT 143.070 154.440 144.470 154.720 ;
        RECT 153.990 154.440 156.790 154.720 ;
        RECT 163.790 154.440 164.910 154.720 ;
        RECT 167.710 154.440 168.270 154.720 ;
        RECT 143.350 154.160 145.030 154.440 ;
        RECT 153.150 154.160 155.950 154.440 ;
        RECT 163.230 154.160 164.350 154.440 ;
        RECT 167.430 154.160 167.990 154.440 ;
        RECT 173.310 154.160 174.150 155.000 ;
        RECT 175.830 154.720 176.670 155.000 ;
        RECT 192.070 154.720 193.190 155.000 ;
        RECT 193.750 154.720 194.590 155.000 ;
        RECT 204.390 154.720 206.070 155.000 ;
        RECT 207.050 154.860 207.470 155.000 ;
        RECT 176.110 154.440 176.950 154.720 ;
        RECT 191.230 154.440 192.350 154.720 ;
        RECT 194.030 154.440 194.870 154.720 ;
        RECT 204.110 154.440 205.790 154.720 ;
        RECT 176.670 154.160 177.230 154.440 ;
        RECT 190.390 154.160 191.790 154.440 ;
        RECT 194.310 154.160 195.150 154.440 ;
        RECT 203.830 154.160 205.510 154.440 ;
        RECT 143.630 153.880 145.310 154.160 ;
        RECT 152.590 153.880 155.390 154.160 ;
        RECT 162.670 153.880 163.790 154.160 ;
        RECT 167.150 153.880 167.990 154.160 ;
        RECT 173.590 153.880 174.150 154.160 ;
        RECT 176.950 153.880 177.790 154.160 ;
        RECT 189.550 153.880 190.950 154.160 ;
        RECT 194.870 153.880 195.430 154.160 ;
        RECT 203.550 153.880 205.230 154.160 ;
        RECT 144.190 153.600 145.870 153.880 ;
        RECT 151.750 153.600 154.830 153.880 ;
        RECT 162.110 153.600 163.230 153.880 ;
        RECT 167.150 153.600 167.710 153.880 ;
        RECT 173.590 153.600 174.430 153.880 ;
        RECT 177.510 153.600 178.070 153.880 ;
        RECT 188.990 153.600 190.110 153.880 ;
        RECT 195.150 153.600 195.710 153.880 ;
        RECT 203.270 153.600 204.950 153.880 ;
        RECT 207.190 153.600 207.470 154.860 ;
        RECT 144.470 153.320 146.150 153.600 ;
        RECT 151.190 153.320 154.270 153.600 ;
        RECT 161.550 153.320 162.670 153.600 ;
        RECT 173.870 153.320 174.430 153.600 ;
        RECT 177.790 153.320 178.630 153.600 ;
        RECT 188.150 153.320 189.270 153.600 ;
        RECT 195.430 153.320 195.990 153.600 ;
        RECT 202.990 153.320 204.670 153.600 ;
        RECT 145.030 153.040 146.430 153.320 ;
        RECT 150.350 153.040 153.710 153.320 ;
        RECT 161.270 153.040 162.110 153.320 ;
        RECT 173.870 153.040 174.710 153.320 ;
        RECT 178.070 153.040 178.910 153.320 ;
        RECT 187.310 153.040 188.710 153.320 ;
        RECT 195.710 153.040 196.270 153.320 ;
        RECT 202.710 153.040 204.390 153.320 ;
        RECT 145.310 152.760 146.990 153.040 ;
        RECT 149.790 152.760 153.150 153.040 ;
        RECT 160.710 152.760 161.830 153.040 ;
        RECT 174.150 152.760 174.710 153.040 ;
        RECT 178.630 152.760 179.190 153.040 ;
        RECT 186.470 152.760 187.870 153.040 ;
        RECT 195.990 152.760 196.270 153.040 ;
        RECT 201.590 152.760 204.110 153.040 ;
        RECT 145.590 152.480 147.270 152.760 ;
        RECT 148.950 152.480 152.590 152.760 ;
        RECT 160.150 152.480 161.270 152.760 ;
        RECT 174.430 152.480 174.990 152.760 ;
        RECT 178.910 152.480 179.750 152.760 ;
        RECT 185.910 152.480 187.030 152.760 ;
        RECT 201.310 152.620 201.730 152.760 ;
        RECT 145.870 152.200 147.550 152.480 ;
        RECT 148.390 152.200 152.030 152.480 ;
        RECT 159.590 152.200 160.710 152.480 ;
        RECT 174.430 152.200 175.270 152.480 ;
        RECT 179.470 152.200 180.030 152.480 ;
        RECT 185.070 152.200 186.190 152.480 ;
        RECT 146.430 151.920 151.190 152.200 ;
        RECT 159.030 151.920 160.150 152.200 ;
        RECT 174.710 151.920 175.550 152.200 ;
        RECT 179.750 151.920 180.590 152.200 ;
        RECT 184.230 151.920 185.630 152.200 ;
        RECT 146.710 151.640 150.630 151.920 ;
        RECT 158.470 151.640 159.590 151.920 ;
        RECT 164.910 151.640 165.470 151.920 ;
        RECT 174.990 151.640 175.830 151.920 ;
        RECT 180.030 151.640 180.870 151.920 ;
        RECT 183.390 151.640 184.790 151.920 ;
        RECT 146.990 151.360 150.070 151.640 ;
        RECT 157.910 151.360 159.030 151.640 ;
        RECT 165.190 151.360 165.750 151.640 ;
        RECT 175.270 151.360 176.110 151.640 ;
        RECT 180.590 151.360 181.430 151.640 ;
        RECT 182.830 151.360 183.950 151.640 ;
        RECT 147.270 151.080 149.510 151.360 ;
        RECT 157.350 151.080 158.470 151.360 ;
        RECT 164.070 151.080 164.910 151.360 ;
        RECT 165.470 151.080 166.030 151.360 ;
        RECT 175.550 151.080 176.390 151.360 ;
        RECT 180.870 151.080 183.390 151.360 ;
        RECT 147.830 150.800 149.230 151.080 ;
        RECT 157.070 150.800 157.910 151.080 ;
        RECT 163.510 150.800 164.350 151.080 ;
        RECT 165.750 150.800 166.310 151.080 ;
        RECT 176.110 150.800 176.670 151.080 ;
        RECT 148.110 150.520 149.790 150.800 ;
        RECT 156.510 150.520 157.350 150.800 ;
        RECT 162.950 150.520 164.070 150.800 ;
        RECT 166.030 150.520 166.590 150.800 ;
        RECT 176.390 150.520 176.950 150.800 ;
        RECT 180.310 150.520 181.150 150.800 ;
        RECT 148.390 150.240 150.070 150.520 ;
        RECT 155.950 150.240 156.790 150.520 ;
        RECT 162.390 150.240 163.790 150.520 ;
        RECT 166.310 150.240 166.870 150.520 ;
        RECT 176.670 150.240 177.230 150.520 ;
        RECT 179.470 150.240 182.270 150.520 ;
        RECT 148.390 149.960 150.350 150.240 ;
        RECT 155.390 149.960 156.230 150.240 ;
        RECT 159.870 149.960 160.150 150.240 ;
        RECT 162.110 149.960 164.070 150.240 ;
        RECT 166.590 149.960 167.150 150.240 ;
        RECT 178.910 149.960 182.830 150.240 ;
        RECT 148.390 149.680 150.630 149.960 ;
        RECT 154.830 149.680 155.670 149.960 ;
        RECT 159.030 149.820 160.430 149.960 ;
        RECT 159.030 149.680 159.870 149.820 ;
        RECT 160.150 149.680 160.430 149.820 ;
        RECT 162.110 149.680 164.350 149.960 ;
        RECT 166.870 149.680 167.430 149.960 ;
        RECT 178.070 149.680 183.390 149.960 ;
        RECT 148.390 149.400 150.910 149.680 ;
        RECT 154.270 149.400 155.110 149.680 ;
        RECT 158.470 149.400 159.310 149.680 ;
        RECT 160.150 149.400 160.710 149.680 ;
        RECT 162.390 149.400 164.630 149.680 ;
        RECT 167.150 149.400 167.710 149.680 ;
        RECT 177.510 149.400 183.950 149.680 ;
        RECT 148.110 149.120 151.190 149.400 ;
        RECT 153.710 149.120 154.550 149.400 ;
        RECT 157.910 149.260 158.610 149.400 ;
        RECT 157.910 149.120 158.470 149.260 ;
        RECT 160.430 149.120 160.710 149.400 ;
        RECT 162.670 149.120 164.910 149.400 ;
        RECT 167.430 149.120 167.990 149.400 ;
        RECT 176.670 149.120 184.230 149.400 ;
        RECT 148.110 148.840 151.750 149.120 ;
        RECT 153.150 148.840 153.990 149.120 ;
        RECT 157.350 148.980 158.050 149.120 ;
        RECT 160.570 148.980 160.990 149.120 ;
        RECT 157.350 148.840 157.910 148.980 ;
        RECT 160.710 148.840 160.990 148.980 ;
        RECT 162.670 148.840 165.190 149.120 ;
        RECT 167.710 148.840 168.270 149.120 ;
        RECT 176.110 148.840 178.350 149.120 ;
        RECT 178.910 148.840 184.510 149.120 ;
        RECT 147.830 148.560 152.030 148.840 ;
        RECT 152.870 148.560 153.430 148.840 ;
        RECT 156.790 148.700 157.490 148.840 ;
        RECT 160.850 148.700 161.270 148.840 ;
        RECT 156.790 148.560 157.350 148.700 ;
        RECT 160.990 148.560 161.270 148.700 ;
        RECT 162.950 148.560 165.470 148.840 ;
        RECT 167.990 148.560 168.550 148.840 ;
        RECT 175.550 148.560 177.790 148.840 ;
        RECT 179.190 148.560 185.070 148.840 ;
        RECT 137.190 148.280 143.350 148.560 ;
        RECT 147.830 148.280 152.310 148.560 ;
        RECT 156.790 148.280 157.070 148.560 ;
        RECT 160.990 148.280 161.550 148.560 ;
        RECT 163.230 148.280 165.470 148.560 ;
        RECT 168.270 148.280 168.830 148.560 ;
        RECT 174.710 148.280 177.230 148.560 ;
        RECT 179.190 148.280 185.350 148.560 ;
        RECT 201.310 148.280 201.590 152.620 ;
        RECT 202.990 152.480 203.830 152.760 ;
        RECT 203.270 152.200 203.550 152.480 ;
        RECT 202.430 151.360 203.270 151.640 ;
        RECT 202.430 151.080 202.710 151.360 ;
        RECT 203.130 151.220 203.550 151.360 ;
        RECT 203.270 151.080 203.550 151.220 ;
        RECT 207.190 151.080 207.470 151.920 ;
        RECT 203.270 150.800 203.830 151.080 ;
        RECT 203.550 150.520 203.830 150.800 ;
        RECT 206.910 150.940 207.330 151.080 ;
        RECT 206.910 150.520 207.190 150.940 ;
        RECT 203.690 150.380 204.110 150.520 ;
        RECT 203.830 150.240 204.110 150.380 ;
        RECT 206.630 150.380 207.050 150.520 ;
        RECT 206.630 150.240 206.910 150.380 ;
        RECT 203.970 150.100 204.390 150.240 ;
        RECT 204.110 149.960 204.390 150.100 ;
        RECT 206.070 150.100 206.770 150.240 ;
        RECT 206.070 149.960 206.630 150.100 ;
        RECT 204.250 149.820 204.950 149.960 ;
        RECT 204.390 149.680 204.950 149.820 ;
        RECT 205.510 149.680 206.350 149.960 ;
        RECT 135.510 148.000 144.750 148.280 ;
        RECT 147.550 148.000 152.590 148.280 ;
        RECT 156.510 148.140 156.930 148.280 ;
        RECT 134.670 147.720 137.470 148.000 ;
        RECT 143.070 147.720 145.590 148.000 ;
        RECT 147.550 147.720 150.910 148.000 ;
        RECT 151.190 147.720 152.870 148.000 ;
        RECT 133.550 147.440 136.070 147.720 ;
        RECT 144.470 147.440 146.430 147.720 ;
        RECT 147.270 147.440 150.630 147.720 ;
        RECT 151.470 147.440 153.150 147.720 ;
        RECT 156.510 147.440 156.790 148.140 ;
        RECT 160.710 148.000 161.270 148.280 ;
        RECT 163.510 148.000 165.750 148.280 ;
        RECT 168.550 148.000 169.110 148.280 ;
        RECT 174.150 148.000 176.390 148.280 ;
        RECT 179.190 148.000 185.910 148.280 ;
        RECT 160.150 147.860 160.850 148.000 ;
        RECT 160.150 147.720 160.710 147.860 ;
        RECT 163.790 147.720 166.030 148.000 ;
        RECT 168.830 147.720 169.390 148.000 ;
        RECT 173.590 147.720 175.830 148.000 ;
        RECT 178.070 147.720 186.190 148.000 ;
        RECT 159.590 147.580 160.290 147.720 ;
        RECT 159.590 147.440 160.150 147.580 ;
        RECT 164.070 147.440 166.310 147.720 ;
        RECT 169.110 147.440 169.670 147.720 ;
        RECT 173.590 147.440 175.270 147.720 ;
        RECT 177.230 147.440 179.190 147.720 ;
        RECT 179.750 147.440 186.470 147.720 ;
        RECT 132.990 147.160 134.950 147.440 ;
        RECT 145.310 147.160 150.630 147.440 ;
        RECT 151.750 147.160 153.430 147.440 ;
        RECT 156.510 147.160 157.070 147.440 ;
        RECT 159.030 147.300 159.730 147.440 ;
        RECT 159.030 147.160 159.590 147.300 ;
        RECT 164.350 147.160 166.590 147.440 ;
        RECT 169.390 147.160 169.950 147.440 ;
        RECT 132.150 146.880 134.110 147.160 ;
        RECT 146.150 146.880 150.350 147.160 ;
        RECT 152.310 146.880 153.710 147.160 ;
        RECT 156.790 146.880 157.070 147.160 ;
        RECT 158.190 147.020 159.170 147.160 ;
        RECT 158.190 146.880 159.030 147.020 ;
        RECT 164.630 146.880 166.870 147.160 ;
        RECT 169.670 146.880 170.230 147.160 ;
        RECT 173.310 146.880 174.430 147.440 ;
        RECT 176.390 147.160 177.510 147.440 ;
        RECT 177.790 147.160 178.350 147.440 ;
        RECT 179.750 147.160 187.030 147.440 ;
        RECT 175.550 146.880 176.950 147.160 ;
        RECT 178.630 146.880 179.190 147.160 ;
        RECT 179.750 146.880 187.310 147.160 ;
        RECT 131.590 146.600 133.270 146.880 ;
        RECT 146.710 146.600 150.350 146.880 ;
        RECT 152.590 146.600 153.990 146.880 ;
        RECT 156.790 146.600 157.350 146.880 ;
        RECT 157.630 146.600 158.470 146.880 ;
        RECT 164.910 146.600 167.150 146.880 ;
        RECT 169.950 146.600 170.510 146.880 ;
        RECT 173.310 146.600 174.150 146.880 ;
        RECT 174.990 146.600 176.390 146.880 ;
        RECT 178.070 146.740 178.770 146.880 ;
        RECT 178.070 146.600 178.630 146.740 ;
        RECT 179.750 146.600 186.190 146.880 ;
        RECT 187.030 146.600 187.870 146.880 ;
        RECT 201.590 146.600 201.870 148.000 ;
        RECT 202.430 147.160 202.710 149.680 ;
        RECT 209.150 148.000 211.110 148.280 ;
        RECT 208.870 147.860 209.290 148.000 ;
        RECT 208.870 147.720 209.150 147.860 ;
        RECT 210.830 147.720 211.390 148.000 ;
        RECT 219.790 147.720 222.590 148.000 ;
        RECT 208.590 147.580 209.010 147.720 ;
        RECT 208.590 147.160 208.870 147.580 ;
        RECT 211.110 147.440 211.670 147.720 ;
        RECT 202.570 147.020 202.990 147.160 ;
        RECT 130.750 146.320 132.430 146.600 ;
        RECT 130.190 146.040 131.870 146.320 ;
        RECT 135.790 146.040 142.230 146.320 ;
        RECT 146.710 146.040 150.070 146.600 ;
        RECT 152.870 146.320 154.270 146.600 ;
        RECT 157.070 146.460 157.770 146.600 ;
        RECT 157.070 146.320 157.630 146.460 ;
        RECT 164.910 146.320 167.430 146.600 ;
        RECT 170.230 146.320 170.790 146.600 ;
        RECT 173.310 146.320 175.550 146.600 ;
        RECT 177.230 146.460 178.210 146.600 ;
        RECT 177.230 146.320 178.070 146.460 ;
        RECT 179.190 146.320 185.630 146.600 ;
        RECT 187.310 146.320 188.150 146.600 ;
        RECT 201.730 146.460 202.150 146.600 ;
        RECT 153.150 146.040 154.550 146.320 ;
        RECT 165.190 146.040 167.430 146.320 ;
        RECT 170.510 146.040 171.070 146.320 ;
        RECT 129.630 145.760 131.030 146.040 ;
        RECT 134.670 145.760 143.630 146.040 ;
        RECT 146.430 145.760 149.790 146.040 ;
        RECT 153.430 145.760 154.830 146.040 ;
        RECT 165.470 145.760 167.710 146.040 ;
        RECT 170.790 145.760 171.070 146.040 ;
        RECT 173.310 146.040 174.990 146.320 ;
        RECT 176.390 146.040 177.510 146.320 ;
        RECT 178.630 146.040 179.330 146.320 ;
        RECT 180.310 146.040 184.790 146.320 ;
        RECT 187.870 146.040 188.710 146.320 ;
        RECT 129.070 145.480 130.470 145.760 ;
        RECT 133.550 145.480 137.190 145.760 ;
        RECT 141.950 145.480 144.470 145.760 ;
        RECT 146.430 145.480 150.070 145.760 ;
        RECT 153.710 145.480 155.110 145.760 ;
        RECT 165.750 145.480 167.990 145.760 ;
        RECT 170.930 145.620 171.350 145.760 ;
        RECT 171.070 145.480 171.350 145.620 ;
        RECT 173.310 145.480 174.430 146.040 ;
        RECT 175.550 145.760 176.950 146.040 ;
        RECT 179.190 145.760 180.030 146.040 ;
        RECT 180.310 145.760 184.230 146.040 ;
        RECT 188.430 145.760 188.990 146.040 ;
        RECT 174.710 145.480 176.390 145.760 ;
        RECT 178.350 145.620 179.330 145.760 ;
        RECT 178.350 145.480 179.190 145.620 ;
        RECT 180.310 145.480 183.670 145.760 ;
        RECT 188.850 145.620 189.550 145.760 ;
        RECT 196.830 145.620 197.390 145.760 ;
        RECT 188.990 145.480 189.550 145.620 ;
        RECT 196.690 145.480 197.390 145.620 ;
        RECT 201.870 145.480 202.150 146.460 ;
        RECT 202.710 145.480 202.990 147.020 ;
        RECT 208.310 146.880 208.870 147.160 ;
        RECT 211.390 146.880 211.670 147.440 ;
        RECT 219.790 147.440 222.870 147.720 ;
        RECT 225.390 147.440 226.790 148.000 ;
        RECT 219.790 147.160 223.150 147.440 ;
        RECT 219.790 146.880 220.630 147.160 ;
        RECT 222.030 146.880 223.150 147.160 ;
        RECT 225.110 147.160 226.790 147.440 ;
        RECT 225.110 146.880 225.670 147.160 ;
        RECT 206.910 146.600 208.590 146.880 ;
        RECT 211.530 146.740 211.950 146.880 ;
        RECT 206.630 146.460 207.050 146.600 ;
        RECT 206.630 146.320 206.910 146.460 ;
        RECT 206.350 146.040 206.910 146.320 ;
        RECT 206.350 145.760 206.630 146.040 ;
        RECT 207.470 145.760 208.870 146.040 ;
        RECT 206.070 145.620 206.490 145.760 ;
        RECT 207.190 145.620 207.610 145.760 ;
        RECT 67.680 144.660 79.600 144.920 ;
        RECT 67.680 144.610 75.560 144.660 ;
        RECT 50.230 143.100 66.920 143.360 ;
        RECT 55.160 142.220 57.170 142.710 ;
        RECT 76.830 142.380 79.130 144.150 ;
        RECT 86.740 142.300 88.900 145.460 ;
        RECT 95.780 142.220 98.290 145.470 ;
        RECT 128.510 145.200 129.910 145.480 ;
        RECT 132.710 145.200 135.790 145.480 ;
        RECT 143.350 145.200 144.470 145.480 ;
        RECT 128.230 144.920 129.350 145.200 ;
        RECT 132.150 144.920 134.670 145.200 ;
        RECT 144.190 144.920 144.470 145.200 ;
        RECT 146.150 145.200 150.630 145.480 ;
        RECT 153.990 145.200 155.390 145.480 ;
        RECT 166.030 145.200 168.270 145.480 ;
        RECT 171.210 145.340 171.630 145.480 ;
        RECT 171.350 145.200 171.630 145.340 ;
        RECT 173.590 145.200 175.550 145.480 ;
        RECT 177.510 145.200 178.630 145.480 ;
        RECT 179.750 145.200 182.830 145.480 ;
        RECT 189.270 145.200 189.830 145.480 ;
        RECT 195.990 145.200 196.830 145.480 ;
        RECT 197.110 145.200 197.670 145.480 ;
        RECT 202.010 145.340 202.430 145.480 ;
        RECT 202.850 145.340 203.270 145.480 ;
        RECT 146.150 144.920 149.510 145.200 ;
        RECT 149.790 144.920 150.910 145.200 ;
        RECT 154.270 144.920 155.670 145.200 ;
        RECT 166.310 144.920 168.550 145.200 ;
        RECT 171.350 144.920 171.910 145.200 ;
        RECT 173.590 144.920 174.990 145.200 ;
        RECT 176.950 144.920 178.070 145.200 ;
        RECT 179.190 144.920 179.890 145.200 ;
        RECT 180.590 145.060 181.010 145.200 ;
        RECT 180.590 144.920 180.870 145.060 ;
        RECT 181.150 144.920 182.270 145.200 ;
        RECT 195.430 144.920 196.270 145.200 ;
        RECT 127.670 144.640 128.790 144.920 ;
        RECT 131.310 144.640 133.830 144.920 ;
        RECT 127.110 144.360 128.510 144.640 ;
        RECT 130.750 144.360 132.990 144.640 ;
        RECT 145.870 144.360 149.230 144.920 ;
        RECT 150.350 144.640 151.470 144.920 ;
        RECT 154.550 144.640 155.950 144.920 ;
        RECT 166.590 144.640 168.830 144.920 ;
        RECT 171.630 144.640 172.190 144.920 ;
        RECT 173.590 144.640 174.710 144.920 ;
        RECT 176.110 144.640 177.510 144.920 ;
        RECT 179.750 144.780 180.730 144.920 ;
        RECT 179.750 144.640 180.590 144.780 ;
        RECT 181.150 144.640 181.710 144.920 ;
        RECT 194.870 144.640 196.270 144.920 ;
        RECT 197.390 144.640 197.670 145.200 ;
        RECT 150.630 144.360 151.750 144.640 ;
        RECT 154.830 144.360 156.230 144.640 ;
        RECT 166.870 144.360 169.110 144.640 ;
        RECT 171.910 144.360 172.470 144.640 ;
        RECT 173.870 144.360 174.990 144.640 ;
        RECT 175.270 144.360 176.670 144.640 ;
        RECT 178.910 144.500 179.890 144.640 ;
        RECT 178.910 144.360 179.750 144.500 ;
        RECT 126.830 144.080 127.950 144.360 ;
        RECT 130.470 144.080 132.430 144.360 ;
        RECT 126.830 143.800 128.230 144.080 ;
        RECT 129.910 143.800 131.870 144.080 ;
        RECT 145.590 143.800 148.950 144.360 ;
        RECT 150.910 144.080 152.030 144.360 ;
        RECT 155.110 144.080 156.510 144.360 ;
        RECT 166.870 144.080 169.390 144.360 ;
        RECT 172.190 144.080 172.750 144.360 ;
        RECT 173.870 144.080 176.110 144.360 ;
        RECT 178.070 144.080 179.190 144.360 ;
        RECT 181.430 144.080 181.710 144.640 ;
        RECT 194.310 144.360 196.270 144.640 ;
        RECT 197.530 144.500 197.950 144.640 ;
        RECT 194.030 144.080 196.550 144.360 ;
        RECT 197.670 144.080 197.950 144.500 ;
        RECT 202.150 144.360 202.430 145.340 ;
        RECT 202.290 144.220 202.710 144.360 ;
        RECT 151.470 143.800 152.310 144.080 ;
        RECT 155.390 143.800 156.790 144.080 ;
        RECT 167.150 143.800 169.670 144.080 ;
        RECT 172.470 143.800 173.030 144.080 ;
        RECT 174.150 143.800 175.550 144.080 ;
        RECT 177.510 143.800 178.630 144.080 ;
        RECT 180.030 143.800 180.310 144.080 ;
        RECT 193.470 143.940 194.170 144.080 ;
        RECT 193.470 143.800 194.030 143.940 ;
        RECT 127.390 143.520 131.310 143.800 ;
        RECT 127.950 143.240 131.030 143.520 ;
        RECT 145.310 143.240 148.670 143.800 ;
        RECT 151.750 143.520 152.590 143.800 ;
        RECT 155.670 143.520 157.070 143.800 ;
        RECT 167.430 143.520 169.670 143.800 ;
        RECT 172.750 143.520 173.310 143.800 ;
        RECT 174.430 143.520 175.550 143.800 ;
        RECT 176.670 143.520 178.070 143.800 ;
        RECT 179.750 143.520 181.990 143.800 ;
        RECT 193.190 143.520 193.750 143.800 ;
        RECT 194.590 143.520 196.550 144.080 ;
        RECT 197.810 143.940 198.230 144.080 ;
        RECT 197.950 143.520 198.230 143.940 ;
        RECT 202.430 143.800 202.710 144.220 ;
        RECT 202.990 144.080 203.270 145.340 ;
        RECT 206.070 145.200 206.350 145.620 ;
        RECT 207.190 145.480 207.470 145.620 ;
        RECT 208.590 145.480 209.150 145.760 ;
        RECT 206.910 145.200 207.470 145.480 ;
        RECT 208.870 145.200 209.150 145.480 ;
        RECT 205.790 145.060 206.210 145.200 ;
        RECT 205.790 144.920 206.070 145.060 ;
        RECT 206.910 144.920 207.190 145.200 ;
        RECT 209.010 145.060 209.430 145.200 ;
        RECT 205.510 144.780 205.930 144.920 ;
        RECT 206.630 144.780 207.050 144.920 ;
        RECT 205.510 144.360 205.790 144.780 ;
        RECT 206.630 144.640 206.910 144.780 ;
        RECT 209.150 144.640 209.430 145.060 ;
        RECT 206.350 144.360 206.910 144.640 ;
        RECT 209.290 144.500 209.710 144.640 ;
        RECT 209.430 144.360 209.710 144.500 ;
        RECT 205.230 144.220 205.650 144.360 ;
        RECT 205.230 144.080 205.510 144.220 ;
        RECT 206.350 144.080 206.630 144.360 ;
        RECT 209.430 144.080 209.990 144.360 ;
        RECT 203.130 143.940 203.550 144.080 ;
        RECT 202.150 143.520 202.990 143.800 ;
        RECT 152.030 143.240 152.870 143.520 ;
        RECT 155.950 143.240 157.350 143.520 ;
        RECT 167.710 143.240 169.950 143.520 ;
        RECT 172.190 143.380 172.890 143.520 ;
        RECT 172.190 143.240 172.750 143.380 ;
        RECT 173.030 143.240 173.590 143.520 ;
        RECT 174.430 143.240 177.510 143.520 ;
        RECT 180.590 143.240 182.270 143.520 ;
        RECT 192.910 143.380 193.330 143.520 ;
        RECT 192.910 143.240 193.190 143.380 ;
        RECT 194.590 143.240 196.830 143.520 ;
        RECT 198.090 143.380 198.510 143.520 ;
        RECT 128.510 142.960 133.270 143.240 ;
        RECT 127.950 142.680 136.070 142.960 ;
        RECT 145.030 142.680 148.390 143.240 ;
        RECT 152.310 142.960 153.150 143.240 ;
        RECT 156.230 142.960 157.630 143.240 ;
        RECT 167.990 142.960 170.230 143.240 ;
        RECT 171.630 143.100 172.330 143.240 ;
        RECT 171.630 142.960 172.190 143.100 ;
        RECT 173.310 142.960 176.670 143.240 ;
        RECT 181.710 142.960 182.270 143.240 ;
        RECT 192.630 143.100 193.050 143.240 ;
        RECT 192.630 142.960 192.910 143.100 ;
        RECT 152.590 142.680 153.430 142.960 ;
        RECT 156.510 142.680 157.910 142.960 ;
        RECT 168.270 142.680 170.510 142.960 ;
        RECT 171.070 142.680 171.910 142.960 ;
        RECT 174.990 142.680 176.390 142.960 ;
        RECT 177.510 142.680 177.790 142.960 ;
        RECT 181.710 142.680 182.550 142.960 ;
        RECT 127.670 142.400 137.190 142.680 ;
        RECT 127.390 142.120 133.270 142.400 ;
        RECT 135.230 142.120 138.030 142.400 ;
        RECT 144.750 142.120 148.110 142.680 ;
        RECT 150.630 142.400 150.910 142.680 ;
        RECT 152.870 142.400 153.710 142.680 ;
        RECT 156.790 142.400 158.190 142.680 ;
        RECT 168.550 142.400 171.350 142.680 ;
        RECT 175.270 142.400 176.670 142.680 ;
        RECT 177.650 142.540 178.070 142.680 ;
        RECT 150.630 142.120 151.470 142.400 ;
        RECT 153.150 142.120 153.990 142.400 ;
        RECT 156.790 142.120 158.470 142.400 ;
        RECT 168.830 142.120 170.790 142.400 ;
        RECT 175.550 142.120 176.950 142.400 ;
        RECT 177.790 142.120 178.070 142.540 ;
        RECT 181.990 142.400 182.550 142.680 ;
        RECT 192.350 142.680 192.910 142.960 ;
        RECT 194.870 142.960 196.830 143.240 ;
        RECT 198.230 143.240 198.510 143.380 ;
        RECT 200.470 143.380 202.290 143.520 ;
        RECT 200.470 143.240 202.150 143.380 ;
        RECT 202.430 143.240 202.990 143.520 ;
        RECT 203.270 143.240 203.550 143.940 ;
        RECT 204.950 143.800 205.510 144.080 ;
        RECT 206.070 143.940 206.490 144.080 ;
        RECT 204.950 143.520 205.230 143.800 ;
        RECT 206.070 143.520 206.350 143.940 ;
        RECT 209.710 143.800 210.270 144.080 ;
        RECT 211.670 143.800 211.950 146.740 ;
        RECT 219.510 146.600 220.630 146.880 ;
        RECT 219.510 145.480 220.350 146.600 ;
        RECT 222.310 146.320 223.150 146.880 ;
        RECT 219.230 144.080 220.070 145.480 ;
        RECT 222.030 144.920 222.870 146.320 ;
        RECT 224.830 146.040 225.670 146.880 ;
        RECT 224.550 145.200 225.390 146.040 ;
        RECT 209.990 143.520 210.550 143.800 ;
        RECT 211.390 143.660 211.810 143.800 ;
        RECT 211.390 143.520 211.670 143.660 ;
        RECT 204.670 143.380 205.090 143.520 ;
        RECT 205.790 143.380 206.210 143.520 ;
        RECT 210.410 143.380 211.530 143.520 ;
        RECT 204.670 143.240 204.950 143.380 ;
        RECT 205.790 143.240 206.070 143.380 ;
        RECT 210.550 143.240 211.390 143.380 ;
        RECT 198.230 142.960 200.190 143.240 ;
        RECT 202.710 142.960 203.550 143.240 ;
        RECT 192.350 142.400 192.630 142.680 ;
        RECT 194.870 142.400 197.110 142.960 ;
        RECT 202.990 142.680 203.550 142.960 ;
        RECT 204.390 142.960 204.950 143.240 ;
        RECT 205.510 142.960 206.070 143.240 ;
        RECT 206.630 142.960 207.190 143.240 ;
        RECT 218.950 142.960 219.790 144.080 ;
        RECT 221.750 143.800 222.590 144.920 ;
        RECT 224.270 144.640 225.110 145.200 ;
        RECT 225.950 144.640 226.790 147.160 ;
        RECT 228.750 146.880 230.150 148.000 ;
        RECT 231.830 147.160 232.670 148.000 ;
        RECT 228.470 146.320 230.150 146.880 ;
        RECT 228.470 145.480 229.310 146.320 ;
        RECT 224.270 144.360 224.830 144.640 ;
        RECT 225.950 144.360 226.510 144.640 ;
        RECT 223.990 143.800 224.830 144.360 ;
        RECT 204.390 142.680 207.190 142.960 ;
        RECT 207.470 142.680 207.750 142.960 ;
        RECT 218.670 142.680 219.790 142.960 ;
        RECT 221.470 143.520 222.590 143.800 ;
        RECT 203.270 142.400 203.830 142.680 ;
        RECT 204.110 142.540 204.530 142.680 ;
        RECT 204.110 142.400 204.390 142.540 ;
        RECT 206.070 142.400 206.630 142.680 ;
        RECT 207.610 142.540 208.030 142.680 ;
        RECT 207.750 142.400 208.030 142.540 ;
        RECT 127.110 141.840 132.710 142.120 ;
        RECT 134.390 141.840 138.590 142.120 ;
        RECT 126.830 141.560 132.150 141.840 ;
        RECT 133.830 141.560 138.870 141.840 ;
        RECT 144.470 141.560 147.830 142.120 ;
        RECT 150.910 141.840 151.750 142.120 ;
        RECT 153.430 141.840 154.270 142.120 ;
        RECT 157.070 141.840 158.750 142.120 ;
        RECT 169.110 141.840 170.230 142.120 ;
        RECT 175.830 141.840 176.950 142.120 ;
        RECT 177.930 141.980 178.350 142.120 ;
        RECT 151.190 141.560 152.030 141.840 ;
        RECT 153.710 141.560 154.550 141.840 ;
        RECT 157.350 141.560 159.030 141.840 ;
        RECT 126.550 141.280 131.590 141.560 ;
        RECT 133.270 141.280 139.430 141.560 ;
        RECT 126.270 141.000 131.310 141.280 ;
        RECT 132.710 141.000 137.190 141.280 ;
        RECT 138.590 141.000 139.710 141.280 ;
        RECT 144.190 141.000 147.550 141.560 ;
        RECT 151.470 141.280 152.310 141.560 ;
        RECT 153.990 141.280 154.830 141.560 ;
        RECT 157.630 141.280 159.030 141.560 ;
        RECT 176.110 141.280 177.230 141.840 ;
        RECT 178.070 141.560 178.350 141.980 ;
        RECT 181.990 141.840 182.830 142.400 ;
        RECT 182.270 141.560 182.830 141.840 ;
        RECT 192.070 142.260 192.490 142.400 ;
        RECT 192.070 141.560 192.350 142.260 ;
        RECT 195.150 141.840 197.390 142.400 ;
        RECT 203.270 142.260 204.250 142.400 ;
        RECT 205.790 142.260 206.210 142.400 ;
        RECT 207.890 142.260 208.310 142.400 ;
        RECT 203.270 142.120 204.110 142.260 ;
        RECT 205.790 142.120 206.070 142.260 ;
        RECT 208.030 142.120 208.310 142.260 ;
        RECT 203.550 141.840 204.110 142.120 ;
        RECT 205.510 141.980 205.930 142.120 ;
        RECT 178.210 141.420 178.630 141.560 ;
        RECT 151.750 141.000 152.590 141.280 ;
        RECT 154.270 141.000 155.110 141.280 ;
        RECT 157.910 141.000 159.310 141.280 ;
        RECT 175.830 141.000 177.510 141.280 ;
        RECT 178.350 141.000 178.630 141.420 ;
        RECT 182.270 141.280 183.110 141.560 ;
        RECT 195.430 141.280 197.670 141.840 ;
        RECT 205.510 141.560 205.790 141.980 ;
        RECT 207.470 141.840 212.230 142.120 ;
        RECT 207.190 141.560 210.830 141.840 ;
        RECT 212.090 141.700 212.510 141.840 ;
        RECT 212.230 141.560 212.510 141.700 ;
        RECT 218.670 141.560 219.510 142.680 ;
        RECT 221.470 142.400 222.310 143.520 ;
        RECT 223.710 142.960 224.550 143.800 ;
        RECT 221.190 142.120 222.310 142.400 ;
        RECT 223.430 142.680 224.270 142.960 ;
        RECT 225.670 142.680 226.510 144.360 ;
        RECT 228.190 144.080 229.030 145.480 ;
        RECT 227.910 142.960 228.750 144.080 ;
        RECT 223.430 142.120 226.510 142.680 ;
        RECT 205.230 141.420 205.650 141.560 ;
        RECT 125.990 140.720 130.750 141.000 ;
        RECT 132.150 140.720 136.070 141.000 ;
        RECT 139.150 140.720 139.990 141.000 ;
        RECT 125.710 140.440 130.470 140.720 ;
        RECT 131.590 140.440 135.230 140.720 ;
        RECT 139.430 140.440 139.990 140.720 ;
        RECT 143.910 140.440 147.270 141.000 ;
        RECT 152.030 140.720 152.870 141.000 ;
        RECT 154.550 140.720 155.390 141.000 ;
        RECT 158.190 140.720 159.590 141.000 ;
        RECT 175.270 140.860 175.970 141.000 ;
        RECT 175.270 140.720 175.830 140.860 ;
        RECT 176.670 140.720 177.510 141.000 ;
        RECT 178.490 140.860 178.910 141.000 ;
        RECT 152.310 140.440 153.150 140.720 ;
        RECT 154.830 140.440 155.390 140.720 ;
        RECT 158.470 140.440 159.870 140.720 ;
        RECT 174.430 140.580 175.410 140.720 ;
        RECT 174.430 140.440 175.270 140.580 ;
        RECT 176.670 140.440 177.790 140.720 ;
        RECT 125.430 140.160 130.190 140.440 ;
        RECT 131.310 140.160 134.390 140.440 ;
        RECT 139.430 140.160 140.270 140.440 ;
        RECT 143.910 140.160 146.990 140.440 ;
        RECT 152.590 140.160 153.430 140.440 ;
        RECT 154.830 140.160 155.670 140.440 ;
        RECT 158.750 140.160 160.150 140.440 ;
        RECT 173.870 140.160 174.710 140.440 ;
        RECT 176.950 140.160 177.790 140.440 ;
        RECT 178.630 140.440 178.910 140.860 ;
        RECT 182.550 140.720 183.110 141.280 ;
        RECT 182.550 140.440 183.390 140.720 ;
        RECT 192.070 140.440 192.350 141.280 ;
        RECT 195.710 140.720 197.950 141.280 ;
        RECT 195.990 140.440 198.230 140.720 ;
        RECT 198.790 140.440 199.070 140.720 ;
        RECT 205.230 140.440 205.510 141.420 ;
        RECT 206.910 141.280 210.830 141.560 ;
        RECT 212.370 141.420 212.790 141.560 ;
        RECT 178.630 140.160 179.190 140.440 ;
        RECT 125.430 139.880 129.630 140.160 ;
        RECT 131.030 139.880 133.830 140.160 ;
        RECT 139.710 139.880 140.550 140.160 ;
        RECT 125.150 139.600 129.350 139.880 ;
        RECT 130.470 139.600 133.270 139.880 ;
        RECT 139.990 139.600 140.550 139.880 ;
        RECT 143.630 139.880 146.990 140.160 ;
        RECT 152.870 139.880 153.430 140.160 ;
        RECT 155.110 139.880 155.950 140.160 ;
        RECT 159.030 139.880 160.430 140.160 ;
        RECT 173.310 139.880 174.150 140.160 ;
        RECT 143.630 139.600 146.710 139.880 ;
        RECT 152.870 139.600 153.710 139.880 ;
        RECT 155.390 139.600 156.230 139.880 ;
        RECT 124.870 139.320 129.070 139.600 ;
        RECT 130.190 139.320 132.990 139.600 ;
        RECT 139.990 139.320 140.830 139.600 ;
        RECT 124.590 139.040 128.790 139.320 ;
        RECT 129.910 139.040 132.430 139.320 ;
        RECT 124.590 138.760 128.510 139.040 ;
        RECT 129.630 138.760 132.150 139.040 ;
        RECT 124.310 138.480 128.230 138.760 ;
        RECT 129.350 138.480 131.590 138.760 ;
        RECT 140.270 138.480 140.830 139.320 ;
        RECT 143.350 139.040 146.710 139.600 ;
        RECT 153.150 139.320 153.990 139.600 ;
        RECT 155.670 139.320 156.230 139.600 ;
        RECT 159.310 139.600 160.710 139.880 ;
        RECT 172.470 139.600 173.590 139.880 ;
        RECT 177.230 139.600 178.070 140.160 ;
        RECT 178.910 139.880 179.190 140.160 ;
        RECT 182.830 139.880 183.390 140.440 ;
        RECT 192.210 140.300 192.630 140.440 ;
        RECT 192.350 139.880 192.630 140.300 ;
        RECT 195.990 140.160 198.510 140.440 ;
        RECT 205.370 140.300 205.790 140.440 ;
        RECT 196.270 139.880 197.950 140.160 ;
        RECT 205.510 139.880 205.790 140.300 ;
        RECT 206.630 140.160 210.550 141.280 ;
        RECT 212.510 140.160 212.790 141.420 ;
        RECT 218.390 140.440 219.230 141.560 ;
        RECT 221.190 141.000 222.030 142.120 ;
        RECT 223.150 141.840 226.510 142.120 ;
        RECT 223.150 141.280 223.990 141.840 ;
        RECT 220.910 140.720 221.750 141.000 ;
        RECT 222.870 140.720 223.710 141.280 ;
        RECT 220.630 140.440 221.750 140.720 ;
        RECT 222.590 140.440 223.710 140.720 ;
        RECT 225.670 140.440 226.510 141.840 ;
        RECT 227.630 142.680 228.750 142.960 ;
        RECT 227.630 141.560 228.470 142.680 ;
        RECT 218.390 140.160 221.470 140.440 ;
        RECT 206.910 139.880 210.830 140.160 ;
        RECT 212.230 140.020 212.650 140.160 ;
        RECT 212.230 139.880 212.510 140.020 ;
        RECT 178.910 139.600 179.470 139.880 ;
        RECT 159.310 139.320 160.990 139.600 ;
        RECT 171.910 139.320 173.030 139.600 ;
        RECT 177.510 139.320 178.350 139.600 ;
        RECT 153.430 139.040 154.270 139.320 ;
        RECT 155.670 139.040 156.510 139.320 ;
        RECT 159.590 139.040 161.270 139.320 ;
        RECT 171.070 139.040 172.470 139.320 ;
        RECT 177.230 139.040 178.350 139.320 ;
        RECT 179.190 139.040 179.470 139.600 ;
        RECT 183.110 139.040 183.670 139.880 ;
        RECT 192.490 139.740 192.910 139.880 ;
        RECT 192.630 139.600 192.910 139.740 ;
        RECT 196.270 139.600 197.390 139.880 ;
        RECT 205.510 139.600 206.070 139.880 ;
        RECT 207.190 139.600 211.110 139.880 ;
        RECT 211.950 139.600 212.510 139.880 ;
        RECT 218.110 139.880 221.190 140.160 ;
        RECT 222.590 139.880 223.430 140.440 ;
        RECT 225.390 139.880 226.510 140.440 ;
        RECT 227.350 140.160 228.190 141.560 ;
        RECT 229.590 141.280 230.150 146.320 ;
        RECT 231.550 146.880 232.670 147.160 ;
        RECT 234.070 146.880 234.910 148.000 ;
        RECT 236.310 147.720 239.110 148.000 ;
        RECT 236.310 147.160 238.830 147.720 ;
        RECT 236.310 146.880 237.150 147.160 ;
        RECT 239.950 146.880 240.790 148.000 ;
        RECT 244.710 147.160 247.790 148.000 ;
        RECT 248.910 147.720 251.710 148.000 ;
        RECT 248.910 147.160 251.430 147.720 ;
        RECT 252.270 147.160 255.350 148.000 ;
        RECT 246.670 146.880 247.510 147.160 ;
        RECT 248.910 146.880 249.750 147.160 ;
        RECT 254.230 146.880 255.070 147.160 ;
        RECT 256.190 146.880 257.590 148.000 ;
        RECT 259.270 147.160 260.110 148.000 ;
        RECT 231.550 145.760 232.390 146.880 ;
        RECT 231.270 145.480 232.390 145.760 ;
        RECT 233.790 146.600 234.910 146.880 ;
        RECT 236.030 146.600 237.150 146.880 ;
        RECT 239.670 146.600 240.790 146.880 ;
        RECT 233.790 145.480 234.630 146.600 ;
        RECT 236.030 145.480 236.870 146.600 ;
        RECT 239.670 145.480 240.510 146.600 ;
        RECT 246.390 146.320 247.230 146.880 ;
        RECT 248.630 146.600 249.750 146.880 ;
        RECT 246.110 145.760 246.950 146.320 ;
        RECT 231.270 144.360 232.110 145.480 ;
        RECT 230.990 143.240 231.830 144.360 ;
        RECT 233.510 144.080 234.350 145.480 ;
        RECT 235.750 144.360 236.590 145.480 ;
        RECT 235.750 144.080 237.990 144.360 ;
        RECT 239.390 144.080 240.230 145.480 ;
        RECT 245.830 145.200 246.670 145.760 ;
        RECT 248.630 145.480 249.470 146.600 ;
        RECT 253.950 146.320 254.790 146.880 ;
        RECT 255.910 146.320 257.590 146.880 ;
        RECT 253.670 145.760 254.510 146.320 ;
        RECT 245.550 144.640 246.390 145.200 ;
        RECT 245.270 144.080 246.110 144.640 ;
        RECT 248.350 144.360 249.190 145.480 ;
        RECT 253.390 145.200 254.230 145.760 ;
        RECT 255.910 145.480 256.750 146.320 ;
        RECT 253.110 144.640 253.950 145.200 ;
        RECT 248.350 144.080 250.590 144.360 ;
        RECT 252.830 144.080 253.670 144.640 ;
        RECT 255.630 144.080 256.470 145.480 ;
        RECT 230.710 142.960 231.830 143.240 ;
        RECT 233.230 142.960 234.070 144.080 ;
        RECT 235.470 143.520 237.990 144.080 ;
        RECT 235.470 142.960 236.310 143.520 ;
        RECT 239.110 142.960 239.950 144.080 ;
        RECT 244.990 143.520 245.830 144.080 ;
        RECT 248.070 143.520 250.590 144.080 ;
        RECT 252.550 143.520 253.390 144.080 ;
        RECT 244.710 142.960 245.550 143.520 ;
        RECT 248.070 142.960 248.910 143.520 ;
        RECT 252.270 142.960 253.110 143.520 ;
        RECT 255.350 142.960 256.190 144.080 ;
        RECT 230.710 141.560 231.550 142.960 ;
        RECT 232.950 142.680 234.070 142.960 ;
        RECT 235.190 142.680 236.310 142.960 ;
        RECT 238.830 142.680 239.950 142.960 ;
        RECT 232.950 141.560 233.790 142.680 ;
        RECT 235.190 141.560 236.030 142.680 ;
        RECT 238.830 141.560 239.670 142.680 ;
        RECT 244.430 142.400 245.270 142.960 ;
        RECT 247.790 142.680 248.910 142.960 ;
        RECT 244.150 141.840 244.990 142.400 ;
        RECT 243.870 141.560 244.710 141.840 ;
        RECT 247.790 141.560 248.630 142.680 ;
        RECT 251.990 142.400 252.830 142.960 ;
        RECT 255.070 142.680 256.190 142.960 ;
        RECT 251.710 141.840 252.550 142.400 ;
        RECT 251.430 141.560 252.270 141.840 ;
        RECT 255.070 141.560 255.910 142.680 ;
        RECT 230.430 141.280 231.270 141.560 ;
        RECT 229.590 140.440 231.270 141.280 ;
        RECT 218.110 139.600 220.910 139.880 ;
        RECT 222.310 139.600 223.150 139.880 ;
        RECT 225.390 139.600 226.230 139.880 ;
        RECT 227.070 139.600 227.910 140.160 ;
        RECT 229.590 139.600 230.990 140.440 ;
        RECT 232.670 140.160 233.510 141.560 ;
        RECT 234.910 140.440 235.750 141.560 ;
        RECT 238.550 140.440 239.390 141.560 ;
        RECT 243.590 141.280 244.710 141.560 ;
        RECT 243.590 141.000 244.430 141.280 ;
        RECT 243.310 140.720 244.430 141.000 ;
        RECT 243.310 140.440 244.150 140.720 ;
        RECT 247.510 140.440 248.350 141.560 ;
        RECT 251.150 141.280 252.270 141.560 ;
        RECT 251.150 141.000 251.990 141.280 ;
        RECT 250.870 140.720 251.990 141.000 ;
        RECT 250.870 140.440 251.710 140.720 ;
        RECT 234.910 140.160 237.430 140.440 ;
        RECT 238.550 140.160 241.070 140.440 ;
        RECT 232.390 139.600 233.230 140.160 ;
        RECT 234.630 139.600 237.430 140.160 ;
        RECT 238.270 139.600 240.790 140.160 ;
        RECT 243.030 139.600 246.110 140.440 ;
        RECT 247.510 140.160 250.030 140.440 ;
        RECT 247.230 139.600 250.030 140.160 ;
        RECT 250.590 139.600 253.670 140.440 ;
        RECT 254.790 140.160 255.630 141.560 ;
        RECT 257.030 141.280 257.590 146.320 ;
        RECT 258.990 146.880 260.110 147.160 ;
        RECT 261.510 146.880 262.350 148.000 ;
        RECT 264.590 147.720 266.550 148.000 ;
        RECT 264.310 147.440 266.830 147.720 ;
        RECT 263.750 147.160 266.830 147.440 ;
        RECT 263.750 146.880 264.870 147.160 ;
        RECT 258.990 145.760 259.830 146.880 ;
        RECT 258.710 145.480 259.830 145.760 ;
        RECT 261.230 146.600 262.350 146.880 ;
        RECT 263.470 146.600 264.590 146.880 ;
        RECT 261.230 145.480 262.070 146.600 ;
        RECT 263.470 145.760 264.310 146.600 ;
        RECT 263.190 145.480 264.310 145.760 ;
        RECT 265.990 146.320 267.110 147.160 ;
        RECT 268.230 146.880 269.070 148.000 ;
        RECT 271.030 147.720 272.150 148.000 ;
        RECT 271.030 147.440 271.870 147.720 ;
        RECT 270.750 147.160 271.590 147.440 ;
        RECT 267.950 146.600 269.070 146.880 ;
        RECT 270.470 146.880 271.590 147.160 ;
        RECT 270.470 146.600 271.310 146.880 ;
        RECT 258.710 144.360 259.550 145.480 ;
        RECT 258.430 143.240 259.270 144.360 ;
        RECT 260.950 144.080 261.790 145.480 ;
        RECT 263.190 144.360 264.030 145.480 ;
        RECT 265.990 145.200 266.830 146.320 ;
        RECT 267.950 145.480 268.790 146.600 ;
        RECT 270.190 146.040 271.030 146.600 ;
        RECT 269.910 145.760 270.750 146.040 ;
        RECT 269.630 145.480 270.750 145.760 ;
        RECT 265.710 144.920 266.550 145.200 ;
        RECT 267.670 144.360 268.510 145.480 ;
        RECT 269.630 145.200 270.470 145.480 ;
        RECT 269.350 144.640 270.190 145.200 ;
        RECT 269.070 144.360 269.910 144.640 ;
        RECT 258.150 142.960 259.270 143.240 ;
        RECT 260.670 142.960 261.510 144.080 ;
        RECT 262.910 142.960 263.750 144.360 ;
        RECT 267.670 144.080 269.630 144.360 ;
        RECT 267.390 143.520 269.630 144.080 ;
        RECT 267.390 142.960 268.230 143.520 ;
        RECT 258.150 141.560 258.990 142.960 ;
        RECT 260.390 142.680 261.510 142.960 ;
        RECT 260.390 141.560 261.230 142.680 ;
        RECT 262.630 141.840 263.470 142.960 ;
        RECT 267.110 142.680 268.230 142.960 ;
        RECT 268.790 142.960 269.630 143.520 ;
        RECT 262.350 141.560 263.470 141.840 ;
        RECT 265.150 142.400 266.270 142.680 ;
        RECT 257.870 141.280 258.710 141.560 ;
        RECT 257.030 140.440 258.710 141.280 ;
        RECT 254.510 139.600 255.350 140.160 ;
        RECT 257.030 139.600 258.430 140.440 ;
        RECT 260.110 140.160 260.950 141.560 ;
        RECT 262.350 140.720 263.190 141.560 ;
        RECT 265.150 141.280 265.990 142.400 ;
        RECT 267.110 141.560 267.950 142.680 ;
        RECT 268.790 142.400 269.910 142.960 ;
        RECT 269.070 141.560 269.910 142.400 ;
        RECT 264.870 141.000 265.990 141.280 ;
        RECT 264.870 140.720 265.710 141.000 ;
        RECT 262.350 140.440 263.470 140.720 ;
        RECT 264.590 140.440 265.710 140.720 ;
        RECT 262.350 140.160 265.430 140.440 ;
        RECT 266.830 140.160 267.670 141.560 ;
        RECT 269.070 141.000 270.190 141.560 ;
        RECT 269.350 140.160 270.190 141.000 ;
        RECT 259.830 139.600 260.670 140.160 ;
        RECT 262.630 139.880 265.150 140.160 ;
        RECT 262.910 139.600 264.870 139.880 ;
        RECT 266.550 139.600 267.390 140.160 ;
        RECT 269.350 139.600 270.470 140.160 ;
        RECT 192.630 139.320 193.190 139.600 ;
        RECT 195.990 139.320 196.830 139.600 ;
        RECT 205.790 139.320 206.350 139.600 ;
        RECT 207.470 139.320 208.030 139.600 ;
        RECT 210.830 139.320 211.110 139.600 ;
        RECT 192.910 139.040 193.470 139.320 ;
        RECT 195.150 139.180 196.130 139.320 ;
        RECT 206.210 139.180 207.610 139.320 ;
        RECT 195.150 139.040 195.990 139.180 ;
        RECT 206.350 139.040 207.470 139.180 ;
        RECT 143.070 138.480 146.430 139.040 ;
        RECT 153.710 138.760 154.550 139.040 ;
        RECT 155.950 138.760 156.790 139.040 ;
        RECT 159.870 138.760 161.270 139.040 ;
        RECT 170.230 138.760 171.910 139.040 ;
        RECT 176.950 138.900 177.370 139.040 ;
        RECT 176.950 138.760 177.230 138.900 ;
        RECT 153.990 138.480 154.830 138.760 ;
        RECT 124.030 137.920 127.950 138.480 ;
        RECT 129.070 138.200 131.310 138.480 ;
        RECT 128.790 137.920 131.030 138.200 ;
        RECT 140.270 137.920 141.110 138.480 ;
        RECT 142.790 137.920 146.150 138.480 ;
        RECT 154.270 138.200 154.830 138.480 ;
        RECT 156.230 138.200 157.070 138.760 ;
        RECT 160.150 138.480 161.550 138.760 ;
        RECT 169.390 138.480 171.350 138.760 ;
        RECT 176.670 138.480 177.230 138.760 ;
        RECT 177.790 138.480 178.630 139.040 ;
        RECT 179.330 138.900 179.750 139.040 ;
        RECT 179.470 138.480 179.750 138.900 ;
        RECT 183.390 138.480 183.950 139.040 ;
        RECT 193.330 138.900 195.430 139.040 ;
        RECT 193.470 138.760 195.430 138.900 ;
        RECT 199.350 138.760 202.150 139.040 ;
        RECT 206.630 138.760 207.190 139.040 ;
        RECT 194.030 138.480 194.870 138.760 ;
        RECT 198.790 138.480 199.630 138.760 ;
        RECT 201.590 138.620 206.770 138.760 ;
        RECT 201.590 138.480 206.630 138.620 ;
        RECT 160.430 138.200 161.830 138.480 ;
        RECT 168.550 138.200 170.510 138.480 ;
        RECT 176.390 138.200 176.950 138.480 ;
        RECT 178.070 138.200 178.910 138.480 ;
        RECT 179.610 138.340 180.030 138.480 ;
        RECT 154.270 137.920 155.110 138.200 ;
        RECT 156.510 137.920 157.350 138.200 ;
        RECT 160.710 137.920 162.110 138.200 ;
        RECT 167.710 137.920 169.950 138.200 ;
        RECT 176.110 137.920 176.670 138.200 ;
        RECT 178.350 137.920 178.910 138.200 ;
        RECT 179.750 137.920 180.030 138.340 ;
        RECT 183.670 138.200 183.950 138.480 ;
        RECT 193.470 138.200 194.310 138.480 ;
        RECT 198.230 138.200 199.070 138.480 ;
        RECT 205.510 138.200 206.630 138.480 ;
        RECT 123.750 137.640 127.670 137.920 ;
        RECT 123.750 137.360 127.390 137.640 ;
        RECT 128.510 137.360 130.750 137.920 ;
        RECT 140.550 137.640 141.110 137.920 ;
        RECT 138.030 137.360 141.110 137.640 ;
        RECT 142.510 137.360 145.870 137.920 ;
        RECT 154.550 137.640 155.390 137.920 ;
        RECT 154.830 137.360 155.390 137.640 ;
        RECT 156.790 137.640 157.350 137.920 ;
        RECT 160.990 137.640 162.390 137.920 ;
        RECT 166.870 137.640 169.390 137.920 ;
        RECT 175.830 137.640 176.390 137.920 ;
        RECT 178.350 137.640 179.190 137.920 ;
        RECT 179.750 137.640 180.310 137.920 ;
        RECT 183.670 137.640 184.230 138.200 ;
        RECT 193.190 137.920 193.750 138.200 ;
        RECT 197.950 137.920 198.510 138.200 ;
        RECT 206.490 138.060 207.190 138.200 ;
        RECT 206.630 137.920 207.190 138.060 ;
        RECT 191.510 137.780 193.330 137.920 ;
        RECT 197.390 137.780 198.090 137.920 ;
        RECT 191.510 137.640 193.190 137.780 ;
        RECT 197.390 137.640 197.950 137.780 ;
        RECT 206.910 137.640 207.470 137.920 ;
        RECT 156.790 137.360 157.630 137.640 ;
        RECT 160.990 137.360 162.670 137.640 ;
        RECT 165.750 137.360 168.550 137.640 ;
        RECT 175.830 137.360 176.110 137.640 ;
        RECT 123.470 137.080 127.110 137.360 ;
        RECT 128.230 137.080 130.470 137.360 ;
        RECT 136.910 137.080 139.150 137.360 ;
        RECT 139.710 137.080 141.110 137.360 ;
        RECT 123.190 136.800 127.110 137.080 ;
        RECT 127.950 136.800 130.470 137.080 ;
        RECT 136.070 136.800 137.470 137.080 ;
        RECT 140.550 136.800 141.110 137.080 ;
        RECT 142.230 137.080 146.710 137.360 ;
        RECT 154.830 137.080 155.670 137.360 ;
        RECT 157.070 137.080 157.910 137.360 ;
        RECT 161.270 137.080 162.670 137.360 ;
        RECT 164.910 137.080 167.710 137.360 ;
        RECT 175.550 137.080 176.110 137.360 ;
        RECT 178.630 137.360 179.190 137.640 ;
        RECT 180.030 137.360 180.310 137.640 ;
        RECT 178.630 137.080 179.470 137.360 ;
        RECT 180.030 137.080 180.590 137.360 ;
        RECT 183.950 137.080 184.510 137.640 ;
        RECT 189.550 137.360 191.790 137.640 ;
        RECT 192.630 137.360 193.190 137.640 ;
        RECT 196.830 137.500 197.530 137.640 ;
        RECT 207.330 137.500 208.030 137.640 ;
        RECT 196.830 137.360 197.390 137.500 ;
        RECT 207.470 137.360 208.030 137.500 ;
        RECT 188.990 137.080 190.390 137.360 ;
        RECT 190.950 137.080 191.230 137.360 ;
        RECT 142.230 136.800 147.550 137.080 ;
        RECT 155.110 136.800 155.950 137.080 ;
        RECT 157.350 136.800 157.910 137.080 ;
        RECT 161.550 136.800 162.950 137.080 ;
        RECT 163.790 136.800 167.150 137.080 ;
        RECT 175.270 136.800 175.830 137.080 ;
        RECT 178.910 136.800 179.470 137.080 ;
        RECT 180.310 136.800 180.590 137.080 ;
        RECT 184.230 136.800 184.510 137.080 ;
        RECT 188.710 136.940 189.130 137.080 ;
        RECT 188.710 136.800 188.990 136.940 ;
        RECT 189.270 136.800 190.390 137.080 ;
        RECT 123.190 136.240 126.830 136.800 ;
        RECT 127.670 136.240 130.470 136.800 ;
        RECT 135.510 136.520 136.630 136.800 ;
        RECT 140.270 136.520 141.110 136.800 ;
        RECT 134.950 136.240 135.790 136.520 ;
        RECT 122.910 135.960 126.550 136.240 ;
        RECT 127.390 135.960 130.470 136.240 ;
        RECT 134.390 135.960 135.230 136.240 ;
        RECT 122.910 135.680 126.270 135.960 ;
        RECT 127.390 135.680 130.750 135.960 ;
        RECT 134.110 135.680 134.950 135.960 ;
        RECT 140.270 135.680 140.830 136.520 ;
        RECT 141.950 136.240 145.310 136.800 ;
        RECT 146.150 136.520 148.390 136.800 ;
        RECT 146.990 136.240 148.950 136.520 ;
        RECT 155.390 136.240 156.230 136.800 ;
        RECT 157.350 136.520 158.190 136.800 ;
        RECT 161.830 136.520 166.310 136.800 ;
        RECT 174.990 136.520 175.550 136.800 ;
        RECT 178.910 136.520 179.750 136.800 ;
        RECT 180.310 136.520 180.870 136.800 ;
        RECT 157.630 136.240 158.190 136.520 ;
        RECT 162.110 136.240 165.470 136.520 ;
        RECT 174.710 136.240 175.270 136.520 ;
        RECT 179.190 136.240 179.750 136.520 ;
        RECT 180.590 136.240 180.870 136.520 ;
        RECT 184.230 136.240 184.790 136.800 ;
        RECT 141.670 135.680 145.030 136.240 ;
        RECT 147.830 135.960 150.070 136.240 ;
        RECT 155.670 135.960 156.510 136.240 ;
        RECT 157.630 135.960 158.470 136.240 ;
        RECT 162.110 135.960 164.630 136.240 ;
        RECT 174.430 135.960 174.990 136.240 ;
        RECT 179.190 135.960 180.030 136.240 ;
        RECT 180.590 135.960 181.150 136.240 ;
        RECT 148.670 135.680 150.910 135.960 ;
        RECT 155.950 135.680 156.510 135.960 ;
        RECT 157.910 135.680 158.470 135.960 ;
        RECT 162.390 135.680 163.790 135.960 ;
        RECT 174.150 135.680 174.710 135.960 ;
        RECT 179.470 135.680 180.030 135.960 ;
        RECT 180.870 135.680 181.150 135.960 ;
        RECT 184.510 135.960 184.790 136.240 ;
        RECT 188.430 136.660 188.850 136.800 ;
        RECT 188.430 135.960 188.710 136.660 ;
        RECT 184.510 135.680 185.070 135.960 ;
        RECT 189.270 135.680 190.110 136.800 ;
        RECT 122.630 135.400 126.270 135.680 ;
        RECT 127.110 135.400 130.750 135.680 ;
        RECT 133.830 135.400 134.390 135.680 ;
        RECT 122.630 134.840 125.990 135.400 ;
        RECT 122.350 134.560 125.990 134.840 ;
        RECT 126.830 135.120 131.030 135.400 ;
        RECT 133.550 135.120 134.110 135.400 ;
        RECT 139.990 135.120 140.830 135.680 ;
        RECT 141.390 135.400 145.030 135.680 ;
        RECT 146.430 135.400 146.710 135.680 ;
        RECT 148.950 135.400 151.750 135.680 ;
        RECT 155.950 135.400 156.790 135.680 ;
        RECT 157.910 135.400 158.750 135.680 ;
        RECT 141.390 135.120 146.710 135.400 ;
        RECT 148.670 135.120 152.590 135.400 ;
        RECT 156.230 135.120 157.070 135.400 ;
        RECT 126.830 134.840 131.310 135.120 ;
        RECT 133.270 134.840 133.830 135.120 ;
        RECT 126.830 134.560 131.870 134.840 ;
        RECT 132.990 134.560 133.550 134.840 ;
        RECT 139.990 134.560 144.470 135.120 ;
        RECT 145.030 134.840 146.990 135.120 ;
        RECT 148.390 134.840 153.710 135.120 ;
        RECT 156.510 134.840 157.070 135.120 ;
        RECT 158.190 135.120 158.750 135.400 ;
        RECT 162.390 135.400 163.230 135.680 ;
        RECT 173.870 135.400 174.430 135.680 ;
        RECT 179.470 135.400 180.310 135.680 ;
        RECT 180.870 135.400 181.430 135.680 ;
        RECT 184.790 135.400 185.070 135.680 ;
        RECT 145.310 134.560 146.990 134.840 ;
        RECT 148.110 134.560 154.550 134.840 ;
        RECT 156.510 134.560 157.350 134.840 ;
        RECT 158.190 134.560 159.030 135.120 ;
        RECT 162.390 134.840 163.510 135.400 ;
        RECT 173.590 135.120 174.150 135.400 ;
        RECT 179.750 135.120 180.310 135.400 ;
        RECT 181.150 135.120 181.430 135.400 ;
        RECT 173.310 134.840 173.870 135.120 ;
        RECT 179.750 134.840 180.590 135.120 ;
        RECT 122.350 134.000 125.710 134.560 ;
        RECT 126.550 134.280 133.270 134.560 ;
        RECT 126.550 134.000 132.990 134.280 ;
        RECT 140.830 134.000 144.190 134.560 ;
        RECT 145.030 134.280 147.270 134.560 ;
        RECT 147.830 134.280 152.310 134.560 ;
        RECT 153.150 134.280 155.950 134.560 ;
        RECT 156.790 134.280 159.030 134.560 ;
        RECT 162.670 134.280 163.790 134.840 ;
        RECT 173.030 134.560 173.590 134.840 ;
        RECT 172.750 134.280 173.310 134.560 ;
        RECT 180.030 134.280 180.590 134.840 ;
        RECT 181.150 134.560 181.710 135.120 ;
        RECT 181.430 134.280 181.710 134.560 ;
        RECT 145.030 134.000 148.950 134.280 ;
        RECT 149.790 134.000 152.590 134.280 ;
        RECT 122.070 133.160 125.430 134.000 ;
        RECT 126.270 133.720 132.710 134.000 ;
        RECT 138.590 133.720 140.270 134.000 ;
        RECT 140.550 133.720 143.910 134.000 ;
        RECT 126.270 133.440 127.950 133.720 ;
        RECT 129.070 133.440 132.710 133.720 ;
        RECT 137.470 133.440 143.910 133.720 ;
        RECT 126.270 133.160 127.670 133.440 ;
        RECT 130.190 133.160 132.430 133.440 ;
        RECT 136.910 133.160 139.150 133.440 ;
        RECT 139.990 133.160 143.630 133.440 ;
        RECT 121.790 132.040 125.150 133.160 ;
        RECT 125.990 132.600 127.670 133.160 ;
        RECT 131.310 132.880 132.150 133.160 ;
        RECT 136.350 132.880 137.750 133.160 ;
        RECT 138.030 132.880 139.150 133.160 ;
        RECT 140.270 132.880 143.630 133.160 ;
        RECT 144.750 132.880 148.670 134.000 ;
        RECT 150.350 133.720 152.590 134.000 ;
        RECT 150.910 133.440 152.590 133.720 ;
        RECT 153.430 134.000 158.470 134.280 ;
        RECT 162.950 134.000 164.070 134.280 ;
        RECT 172.470 134.000 173.030 134.280 ;
        RECT 153.430 133.720 157.910 134.000 ;
        RECT 162.950 133.720 164.350 134.000 ;
        RECT 171.910 133.720 172.750 134.000 ;
        RECT 180.310 133.720 180.870 134.280 ;
        RECT 181.430 134.000 181.990 134.280 ;
        RECT 181.710 133.720 181.990 134.000 ;
        RECT 153.430 133.440 156.790 133.720 ;
        RECT 163.230 133.440 164.350 133.720 ;
        RECT 171.630 133.440 172.470 133.720 ;
        RECT 131.590 132.600 132.150 132.880 ;
        RECT 136.070 132.600 137.190 132.880 ;
        RECT 125.990 132.320 127.390 132.600 ;
        RECT 131.590 132.320 131.870 132.600 ;
        RECT 135.790 132.320 136.630 132.600 ;
        RECT 121.790 131.760 124.870 132.040 ;
        RECT 121.510 130.360 124.870 131.760 ;
        RECT 125.710 131.480 127.390 132.320 ;
        RECT 131.310 132.040 131.870 132.320 ;
        RECT 135.510 132.040 136.350 132.320 ;
        RECT 138.310 132.040 139.150 132.880 ;
        RECT 139.990 132.320 143.350 132.880 ;
        RECT 139.710 132.040 143.350 132.320 ;
        RECT 144.750 132.600 148.390 132.880 ;
        RECT 151.190 132.600 152.870 133.440 ;
        RECT 131.310 131.760 131.590 132.040 ;
        RECT 135.230 131.760 136.070 132.040 ;
        RECT 138.310 131.760 139.430 132.040 ;
        RECT 139.710 131.760 143.630 132.040 ;
        RECT 144.750 131.760 148.670 132.600 ;
        RECT 151.470 131.760 153.150 132.600 ;
        RECT 153.710 132.320 157.070 133.440 ;
        RECT 125.710 130.920 127.110 131.480 ;
        RECT 121.510 127.280 124.590 130.360 ;
        RECT 125.430 128.400 127.110 130.920 ;
        RECT 131.030 131.200 131.590 131.760 ;
        RECT 134.950 131.480 135.790 131.760 ;
        RECT 134.950 131.200 135.510 131.480 ;
        RECT 131.030 130.640 131.310 131.200 ;
        RECT 134.670 130.920 135.510 131.200 ;
        RECT 138.590 131.200 142.790 131.760 ;
        RECT 143.070 131.480 143.910 131.760 ;
        RECT 143.350 131.200 144.190 131.480 ;
        RECT 144.750 131.200 148.950 131.760 ;
        RECT 151.750 131.200 153.150 131.760 ;
        RECT 153.990 132.040 157.070 132.320 ;
        RECT 134.670 130.640 135.230 130.920 ;
        RECT 138.590 130.640 142.510 131.200 ;
        RECT 143.630 130.920 144.190 131.200 ;
        RECT 145.030 130.920 149.510 131.200 ;
        RECT 143.630 130.640 144.470 130.920 ;
        RECT 130.750 129.800 131.310 130.640 ;
        RECT 134.390 130.360 135.230 130.640 ;
        RECT 134.390 130.080 134.950 130.360 ;
        RECT 138.870 130.080 142.230 130.640 ;
        RECT 143.910 130.080 144.470 130.640 ;
        RECT 145.030 130.080 149.790 130.920 ;
        RECT 134.390 129.800 135.790 130.080 ;
        RECT 125.430 128.120 127.670 128.400 ;
        RECT 125.430 127.840 128.510 128.120 ;
        RECT 130.750 127.840 131.030 129.800 ;
        RECT 134.110 129.520 137.750 129.800 ;
        RECT 138.590 129.520 141.950 130.080 ;
        RECT 143.910 129.800 144.750 130.080 ;
        RECT 134.110 129.240 141.670 129.520 ;
        RECT 125.430 127.560 129.630 127.840 ;
        RECT 125.430 127.280 130.470 127.560 ;
        RECT 130.750 127.280 131.310 127.840 ;
        RECT 134.110 127.560 134.670 129.240 ;
        RECT 135.230 128.960 141.670 129.240 ;
        RECT 137.190 128.680 141.670 128.960 ;
        RECT 138.310 128.400 143.350 128.680 ;
        RECT 144.190 128.400 144.750 129.800 ;
        RECT 145.310 129.800 149.790 130.080 ;
        RECT 151.750 129.800 153.430 131.200 ;
        RECT 153.990 130.920 157.350 132.040 ;
        RECT 145.310 129.240 149.510 129.800 ;
        RECT 145.590 128.680 149.510 129.240 ;
        RECT 138.310 127.840 144.750 128.400 ;
        RECT 138.310 127.560 141.110 127.840 ;
        RECT 143.070 127.560 144.750 127.840 ;
        RECT 134.110 127.280 134.950 127.560 ;
        RECT 138.310 127.280 140.830 127.560 ;
        RECT 144.190 127.280 144.750 127.560 ;
        RECT 145.870 127.280 149.230 128.680 ;
        RECT 152.030 127.840 153.430 129.800 ;
        RECT 121.510 126.160 124.870 127.280 ;
        RECT 125.430 127.000 131.310 127.280 ;
        RECT 121.790 125.600 124.870 126.160 ;
        RECT 125.710 126.720 131.310 127.000 ;
        RECT 134.390 126.720 134.950 127.280 ;
        RECT 138.030 127.000 140.830 127.280 ;
        RECT 137.750 126.720 140.830 127.000 ;
        RECT 143.910 127.000 144.750 127.280 ;
        RECT 146.150 127.000 148.950 127.280 ;
        RECT 125.710 126.160 131.590 126.720 ;
        RECT 134.390 126.440 135.230 126.720 ;
        RECT 137.470 126.440 138.870 126.720 ;
        RECT 125.710 125.880 129.910 126.160 ;
        RECT 130.750 125.880 131.590 126.160 ;
        RECT 134.670 126.160 135.230 126.440 ;
        RECT 137.190 126.160 138.590 126.440 ;
        RECT 139.990 126.160 141.110 126.720 ;
        RECT 143.910 126.440 144.470 127.000 ;
        RECT 146.150 126.720 148.670 127.000 ;
        RECT 146.710 126.440 148.390 126.720 ;
        RECT 151.750 126.440 153.430 127.840 ;
        RECT 154.270 126.720 157.350 130.920 ;
        RECT 163.510 130.640 164.350 133.440 ;
        RECT 171.350 133.160 172.190 133.440 ;
        RECT 180.590 133.160 181.150 133.720 ;
        RECT 181.710 133.440 182.270 133.720 ;
        RECT 171.070 132.880 171.910 133.160 ;
        RECT 180.870 132.880 181.150 133.160 ;
        RECT 181.990 133.160 182.270 133.440 ;
        RECT 181.990 132.880 182.550 133.160 ;
        RECT 170.790 132.600 171.630 132.880 ;
        RECT 180.870 132.600 181.430 132.880 ;
        RECT 182.270 132.600 182.550 132.880 ;
        RECT 188.150 132.600 188.430 135.680 ;
        RECT 188.990 134.560 190.110 135.680 ;
        RECT 170.510 132.320 171.350 132.600 ;
        RECT 181.150 132.320 181.430 132.600 ;
        RECT 170.230 132.040 171.070 132.320 ;
        RECT 169.670 131.760 170.790 132.040 ;
        RECT 181.150 131.760 181.710 132.320 ;
        RECT 169.390 131.480 170.510 131.760 ;
        RECT 169.110 131.200 170.230 131.480 ;
        RECT 168.830 130.920 169.670 131.200 ;
        RECT 181.430 130.920 181.710 131.760 ;
        RECT 168.270 130.640 169.390 130.920 ;
        RECT 181.430 130.640 181.990 130.920 ;
        RECT 163.230 130.080 164.350 130.640 ;
        RECT 167.990 130.360 169.110 130.640 ;
        RECT 181.710 130.360 181.990 130.640 ;
        RECT 167.710 130.080 168.830 130.360 ;
        RECT 181.710 130.080 182.270 130.360 ;
        RECT 163.230 129.240 164.070 130.080 ;
        RECT 167.430 129.800 168.270 130.080 ;
        RECT 181.990 129.800 182.550 130.080 ;
        RECT 166.870 129.520 167.990 129.800 ;
        RECT 176.110 129.520 176.390 129.800 ;
        RECT 182.270 129.520 182.830 129.800 ;
        RECT 188.150 129.520 188.430 132.320 ;
        RECT 188.990 129.800 189.830 134.560 ;
        RECT 190.670 134.000 190.950 136.800 ;
        RECT 190.810 133.860 191.230 134.000 ;
        RECT 190.950 133.160 191.230 133.860 ;
        RECT 191.510 133.720 191.790 137.360 ;
        RECT 193.050 137.220 193.470 137.360 ;
        RECT 193.190 137.080 193.470 137.220 ;
        RECT 196.270 137.220 196.970 137.360 ;
        RECT 196.270 137.080 196.830 137.220 ;
        RECT 193.330 136.940 193.750 137.080 ;
        RECT 193.470 136.800 193.750 136.940 ;
        RECT 195.990 136.940 196.410 137.080 ;
        RECT 195.990 136.800 196.270 136.940 ;
        RECT 205.510 136.800 205.790 137.360 ;
        RECT 207.890 137.220 208.590 137.360 ;
        RECT 208.030 137.080 208.590 137.220 ;
        RECT 217.550 137.080 270.750 137.640 ;
        RECT 208.030 136.800 209.150 137.080 ;
        RECT 217.550 136.800 270.470 137.080 ;
        RECT 193.470 136.520 194.030 136.800 ;
        RECT 205.230 136.660 205.650 136.800 ;
        RECT 205.230 136.520 205.510 136.660 ;
        RECT 208.030 136.520 209.430 136.800 ;
        RECT 193.750 136.240 194.030 136.520 ;
        RECT 196.830 136.240 197.390 136.520 ;
        RECT 204.670 136.380 205.370 136.520 ;
        RECT 204.670 136.240 205.230 136.380 ;
        RECT 193.890 136.100 194.310 136.240 ;
        RECT 194.030 135.960 194.310 136.100 ;
        RECT 196.270 136.100 196.970 136.240 ;
        RECT 197.250 136.100 197.950 136.240 ;
        RECT 196.270 135.960 196.830 136.100 ;
        RECT 197.390 135.960 197.950 136.100 ;
        RECT 203.830 135.960 205.230 136.240 ;
        RECT 208.030 136.240 209.990 136.520 ;
        RECT 217.270 136.240 270.190 136.800 ;
        RECT 208.030 135.960 210.270 136.240 ;
        RECT 194.170 135.820 194.590 135.960 ;
        RECT 194.310 134.840 194.590 135.820 ;
        RECT 196.270 135.680 196.550 135.960 ;
        RECT 197.810 135.820 198.230 135.960 ;
        RECT 197.950 135.680 198.230 135.820 ;
        RECT 203.830 135.680 204.110 135.960 ;
        RECT 198.090 135.540 198.790 135.680 ;
        RECT 203.970 135.540 204.390 135.680 ;
        RECT 198.230 135.400 198.790 135.540 ;
        RECT 196.270 135.120 196.550 135.400 ;
        RECT 198.650 135.260 199.070 135.400 ;
        RECT 198.790 135.120 199.070 135.260 ;
        RECT 204.110 135.120 204.390 135.540 ;
        RECT 204.670 135.400 204.950 135.960 ;
        RECT 208.030 135.680 210.830 135.960 ;
        RECT 216.990 135.680 269.910 136.240 ;
        RECT 207.750 135.400 211.110 135.680 ;
        RECT 216.990 135.400 269.630 135.680 ;
        RECT 204.810 135.260 205.510 135.400 ;
        RECT 204.950 135.120 205.510 135.260 ;
        RECT 207.750 135.120 211.390 135.400 ;
        RECT 196.270 134.840 196.830 135.120 ;
        RECT 198.930 134.980 199.350 135.120 ;
        RECT 199.070 134.840 199.350 134.980 ;
        RECT 203.830 134.840 204.390 135.120 ;
        RECT 205.370 134.980 206.350 135.120 ;
        RECT 205.510 134.840 206.350 134.980 ;
        RECT 207.470 134.840 208.030 135.120 ;
        RECT 208.310 134.840 211.670 135.120 ;
        RECT 194.030 133.720 194.590 134.840 ;
        RECT 195.990 134.560 197.110 134.840 ;
        RECT 199.210 134.700 199.630 134.840 ;
        RECT 195.710 134.280 197.390 134.560 ;
        RECT 199.350 134.280 199.630 134.700 ;
        RECT 202.990 134.700 203.970 134.840 ;
        RECT 202.990 134.560 203.830 134.700 ;
        RECT 206.070 134.560 206.910 134.840 ;
        RECT 207.470 134.560 207.750 134.840 ;
        RECT 209.150 134.560 211.670 134.840 ;
        RECT 202.430 134.280 203.270 134.560 ;
        RECT 206.770 134.420 207.610 134.560 ;
        RECT 206.910 134.280 207.470 134.420 ;
        RECT 209.710 134.280 211.670 134.560 ;
        RECT 195.710 134.000 197.950 134.280 ;
        RECT 201.870 134.140 202.570 134.280 ;
        RECT 201.870 134.000 202.430 134.140 ;
        RECT 210.270 134.000 211.670 134.280 ;
        RECT 195.430 133.720 198.510 134.000 ;
        RECT 198.790 133.720 199.350 134.000 ;
        RECT 201.310 133.860 202.010 134.000 ;
        RECT 201.310 133.720 201.870 133.860 ;
        RECT 206.350 133.720 208.310 134.000 ;
        RECT 210.830 133.720 211.390 134.000 ;
        RECT 193.750 133.580 194.170 133.720 ;
        RECT 194.450 133.580 194.870 133.720 ;
        RECT 193.750 133.440 194.030 133.580 ;
        RECT 193.470 133.300 193.890 133.440 ;
        RECT 193.470 133.160 193.750 133.300 ;
        RECT 190.950 132.880 191.510 133.160 ;
        RECT 191.230 132.600 191.510 132.880 ;
        RECT 191.790 132.600 192.070 133.160 ;
        RECT 193.190 132.880 193.750 133.160 ;
        RECT 194.590 133.160 194.870 133.580 ;
        RECT 195.430 133.580 198.930 133.720 ;
        RECT 195.430 133.440 198.790 133.580 ;
        RECT 195.150 133.160 198.230 133.440 ;
        RECT 201.310 133.160 201.590 133.720 ;
        RECT 205.230 133.440 209.990 133.720 ;
        RECT 204.390 133.160 210.830 133.440 ;
        RECT 194.590 132.880 198.230 133.160 ;
        RECT 201.030 133.020 201.450 133.160 ;
        RECT 192.910 132.600 193.470 132.880 ;
        RECT 194.590 132.600 197.950 132.880 ;
        RECT 191.370 132.460 193.050 132.600 ;
        RECT 191.510 132.320 192.910 132.460 ;
        RECT 194.590 132.320 197.670 132.600 ;
        RECT 201.030 132.320 201.310 133.020 ;
        RECT 203.830 132.880 207.190 133.160 ;
        RECT 208.030 132.880 211.670 133.160 ;
        RECT 203.270 132.600 205.790 132.880 ;
        RECT 209.710 132.600 212.510 132.880 ;
        RECT 202.990 132.320 204.950 132.600 ;
        RECT 210.550 132.320 213.070 132.600 ;
        RECT 194.310 132.040 197.670 132.320 ;
        RECT 198.230 132.040 198.510 132.320 ;
        RECT 200.750 132.180 201.170 132.320 ;
        RECT 194.310 131.760 197.390 132.040 ;
        RECT 194.030 131.480 197.390 131.760 ;
        RECT 197.950 131.760 199.070 132.040 ;
        RECT 200.750 131.760 201.030 132.180 ;
        RECT 202.710 132.040 204.110 132.320 ;
        RECT 211.390 132.040 213.630 132.320 ;
        RECT 202.430 131.760 203.830 132.040 ;
        RECT 212.230 131.760 214.190 132.040 ;
        RECT 197.950 131.480 199.630 131.760 ;
        RECT 200.470 131.480 201.030 131.760 ;
        RECT 202.150 131.480 203.270 131.760 ;
        RECT 212.790 131.480 214.750 131.760 ;
        RECT 193.750 131.200 197.110 131.480 ;
        RECT 197.670 131.200 199.910 131.480 ;
        RECT 200.470 131.200 200.750 131.480 ;
        RECT 193.750 130.920 196.830 131.200 ;
        RECT 197.670 130.920 200.750 131.200 ;
        RECT 201.870 130.920 202.990 131.480 ;
        RECT 204.670 131.200 204.950 131.480 ;
        RECT 213.350 131.200 215.310 131.480 ;
        RECT 204.110 131.060 204.810 131.200 ;
        RECT 204.110 130.920 204.670 131.060 ;
        RECT 213.910 130.920 215.590 131.200 ;
        RECT 193.470 130.640 196.830 130.920 ;
        RECT 197.390 130.640 200.470 130.920 ;
        RECT 193.190 130.360 196.550 130.640 ;
        RECT 197.110 130.360 200.470 130.640 ;
        RECT 201.590 130.640 202.710 130.920 ;
        RECT 203.830 130.640 204.390 130.920 ;
        RECT 211.950 130.640 212.510 130.920 ;
        RECT 214.470 130.640 216.150 130.920 ;
        RECT 201.590 130.360 202.430 130.640 ;
        RECT 193.190 130.080 196.270 130.360 ;
        RECT 197.110 130.080 200.190 130.360 ;
        RECT 192.910 129.800 196.270 130.080 ;
        RECT 196.830 129.800 200.190 130.080 ;
        RECT 166.590 129.240 167.710 129.520 ;
        RECT 162.950 128.400 164.070 129.240 ;
        RECT 166.310 128.960 167.150 129.240 ;
        RECT 175.830 128.960 176.670 129.520 ;
        RECT 188.290 129.380 188.710 129.520 ;
        RECT 165.750 128.680 166.870 128.960 ;
        RECT 169.670 128.680 169.950 128.960 ;
        RECT 175.550 128.680 176.390 128.960 ;
        RECT 188.430 128.680 188.710 129.380 ;
        RECT 188.990 128.960 190.110 129.800 ;
        RECT 192.910 129.520 195.990 129.800 ;
        RECT 192.630 129.240 195.990 129.520 ;
        RECT 196.550 129.520 200.190 129.800 ;
        RECT 201.310 130.080 202.430 130.360 ;
        RECT 203.550 130.360 204.110 130.640 ;
        RECT 212.230 130.360 212.790 130.640 ;
        RECT 215.030 130.360 216.710 130.640 ;
        RECT 203.550 130.080 203.830 130.360 ;
        RECT 212.650 130.220 213.350 130.360 ;
        RECT 212.790 130.080 213.350 130.220 ;
        RECT 215.590 130.080 216.990 130.360 ;
        RECT 196.550 129.240 200.470 129.520 ;
        RECT 192.350 128.960 195.710 129.240 ;
        RECT 196.270 128.960 201.030 129.240 ;
        RECT 201.310 128.960 202.150 130.080 ;
        RECT 165.470 128.400 166.310 128.680 ;
        RECT 169.390 128.400 169.950 128.680 ;
        RECT 162.950 128.120 163.790 128.400 ;
        RECT 165.190 128.120 166.030 128.400 ;
        RECT 169.390 128.120 169.670 128.400 ;
        RECT 170.510 128.120 171.350 128.680 ;
        RECT 175.270 128.400 175.830 128.680 ;
        RECT 188.570 128.540 188.990 128.680 ;
        RECT 188.710 128.400 188.990 128.540 ;
        RECT 189.270 128.400 190.110 128.960 ;
        RECT 192.070 128.680 195.430 128.960 ;
        RECT 196.270 128.680 202.150 128.960 ;
        RECT 191.790 128.400 195.430 128.680 ;
        RECT 195.990 128.400 202.150 128.680 ;
        RECT 175.270 128.120 175.550 128.400 ;
        RECT 178.070 128.120 178.630 128.400 ;
        RECT 188.710 128.120 190.110 128.400 ;
        RECT 191.230 128.120 195.150 128.400 ;
        RECT 162.670 127.560 163.790 128.120 ;
        RECT 166.590 127.840 167.430 128.120 ;
        RECT 169.110 127.840 169.670 128.120 ;
        RECT 170.230 127.840 171.070 128.120 ;
        RECT 177.510 127.840 178.910 128.120 ;
        RECT 188.990 127.980 191.370 128.120 ;
        RECT 188.990 127.840 191.230 127.980 ;
        RECT 191.790 127.840 194.870 128.120 ;
        RECT 195.710 127.840 202.150 128.400 ;
        RECT 203.270 129.800 203.830 130.080 ;
        RECT 213.070 129.800 213.910 130.080 ;
        RECT 215.870 129.800 217.550 130.080 ;
        RECT 203.270 128.120 203.550 129.800 ;
        RECT 213.630 129.520 214.190 129.800 ;
        RECT 216.430 129.520 217.830 129.800 ;
        RECT 208.870 129.240 210.270 129.520 ;
        RECT 214.050 129.380 214.750 129.520 ;
        RECT 214.190 129.240 214.750 129.380 ;
        RECT 216.990 129.240 218.390 129.520 ;
        RECT 208.030 128.960 210.830 129.240 ;
        RECT 214.470 128.960 215.030 129.240 ;
        RECT 217.270 128.960 218.670 129.240 ;
        RECT 207.750 128.680 211.390 128.960 ;
        RECT 214.890 128.820 215.590 128.960 ;
        RECT 215.030 128.680 215.590 128.820 ;
        RECT 217.830 128.680 218.950 128.960 ;
        RECT 207.470 128.400 208.590 128.680 ;
        RECT 210.550 128.400 211.670 128.680 ;
        RECT 215.310 128.400 216.150 128.680 ;
        RECT 218.110 128.400 219.510 128.680 ;
        RECT 207.470 128.120 208.310 128.400 ;
        RECT 209.150 128.120 209.990 128.400 ;
        RECT 210.830 128.120 211.670 128.400 ;
        RECT 215.870 128.120 216.430 128.400 ;
        RECT 218.670 128.120 219.790 128.400 ;
        RECT 166.590 127.560 167.710 127.840 ;
        RECT 168.830 127.560 169.390 127.840 ;
        RECT 170.230 127.560 170.510 127.840 ;
        RECT 173.310 127.560 173.870 127.840 ;
        RECT 176.950 127.560 178.910 127.840 ;
        RECT 189.830 127.560 190.390 127.840 ;
        RECT 191.510 127.560 194.870 127.840 ;
        RECT 195.430 127.560 202.430 127.840 ;
        RECT 203.270 127.560 203.830 128.120 ;
        RECT 207.190 127.840 208.030 128.120 ;
        RECT 208.590 127.840 210.550 128.120 ;
        RECT 207.190 127.560 207.750 127.840 ;
        RECT 162.670 127.280 163.510 127.560 ;
        RECT 166.310 127.280 167.430 127.560 ;
        RECT 162.390 126.720 163.510 127.280 ;
        RECT 166.030 127.000 167.430 127.280 ;
        RECT 168.550 127.000 169.110 127.560 ;
        RECT 172.750 127.280 174.150 127.560 ;
        RECT 174.710 127.280 175.550 127.560 ;
        RECT 176.390 127.280 178.630 127.560 ;
        RECT 169.670 127.000 170.230 127.280 ;
        RECT 171.350 127.000 172.190 127.280 ;
        RECT 172.470 127.000 173.870 127.280 ;
        RECT 174.430 127.000 175.550 127.280 ;
        RECT 176.110 127.000 178.350 127.280 ;
        RECT 191.230 127.000 194.590 127.560 ;
        RECT 195.150 127.000 202.430 127.560 ;
        RECT 203.550 127.280 203.830 127.560 ;
        RECT 203.550 127.000 204.110 127.280 ;
        RECT 165.750 126.720 167.430 127.000 ;
        RECT 168.270 126.720 168.830 127.000 ;
        RECT 169.390 126.720 170.230 127.000 ;
        RECT 171.070 126.720 173.870 127.000 ;
        RECT 174.150 126.720 175.270 127.000 ;
        RECT 175.830 126.720 178.350 127.000 ;
        RECT 190.950 126.720 194.310 127.000 ;
        RECT 143.630 126.160 144.470 126.440 ;
        RECT 134.670 125.880 135.510 126.160 ;
        RECT 136.910 125.880 138.310 126.160 ;
        RECT 140.270 125.880 141.110 126.160 ;
        RECT 143.350 125.880 144.190 126.160 ;
        RECT 147.270 125.880 147.830 126.440 ;
        RECT 151.750 126.160 153.150 126.440 ;
        RECT 125.710 125.600 129.070 125.880 ;
        RECT 121.790 124.760 125.150 125.600 ;
        RECT 125.710 125.320 128.790 125.600 ;
        RECT 131.310 125.320 131.870 125.880 ;
        RECT 134.950 125.320 135.790 125.880 ;
        RECT 136.630 125.600 138.030 125.880 ;
        RECT 140.270 125.600 141.390 125.880 ;
        RECT 143.350 125.600 143.910 125.880 ;
        RECT 147.270 125.600 147.550 125.880 ;
        RECT 136.350 125.320 137.750 125.600 ;
        RECT 140.550 125.320 141.390 125.600 ;
        RECT 143.070 125.320 143.910 125.600 ;
        RECT 146.990 125.320 147.550 125.600 ;
        RECT 151.470 125.320 153.150 126.160 ;
        RECT 153.990 125.600 157.350 126.720 ;
        RECT 162.110 126.160 163.230 126.720 ;
        RECT 165.470 126.440 167.430 126.720 ;
        RECT 167.990 126.440 170.230 126.720 ;
        RECT 170.790 126.440 178.350 126.720 ;
        RECT 179.190 126.440 180.030 126.720 ;
        RECT 165.470 126.160 166.030 126.440 ;
        RECT 162.110 125.880 162.950 126.160 ;
        RECT 165.190 125.880 165.750 126.160 ;
        RECT 166.310 125.880 167.150 126.440 ;
        RECT 167.990 126.300 176.110 126.440 ;
        RECT 176.530 126.300 178.070 126.440 ;
        RECT 167.990 126.160 175.970 126.300 ;
        RECT 176.670 126.160 178.070 126.300 ;
        RECT 178.910 126.160 180.030 126.440 ;
        RECT 190.670 126.160 194.030 126.720 ;
        RECT 194.870 126.440 202.710 127.000 ;
        RECT 203.830 126.720 204.110 127.000 ;
        RECT 203.830 126.440 204.390 126.720 ;
        RECT 194.590 126.160 202.710 126.440 ;
        RECT 204.110 126.160 204.390 126.440 ;
        RECT 206.910 126.160 207.750 127.560 ;
        RECT 208.310 127.000 210.830 127.840 ;
        RECT 211.110 127.560 211.950 128.120 ;
        RECT 216.150 127.840 216.990 128.120 ;
        RECT 218.950 127.840 220.350 128.120 ;
        RECT 216.710 127.560 217.270 127.840 ;
        RECT 219.230 127.560 220.630 127.840 ;
        RECT 208.030 126.720 210.830 127.000 ;
        RECT 208.310 126.160 210.830 126.720 ;
        RECT 211.390 126.440 212.230 127.560 ;
        RECT 217.130 127.420 217.830 127.560 ;
        RECT 217.270 127.280 217.830 127.420 ;
        RECT 219.790 127.280 220.910 127.560 ;
        RECT 217.550 127.000 218.390 127.280 ;
        RECT 220.070 127.000 221.190 127.280 ;
        RECT 218.110 126.720 218.670 127.000 ;
        RECT 220.630 126.720 221.750 127.000 ;
        RECT 218.390 126.440 219.230 126.720 ;
        RECT 220.910 126.440 222.030 126.720 ;
        RECT 211.390 126.160 211.950 126.440 ;
        RECT 218.950 126.160 219.510 126.440 ;
        RECT 221.190 126.160 222.310 126.440 ;
        RECT 167.710 125.880 168.550 126.160 ;
        RECT 168.830 125.880 175.830 126.160 ;
        RECT 176.390 125.880 179.470 126.160 ;
        RECT 190.390 125.880 193.750 126.160 ;
        RECT 161.830 125.600 162.950 125.880 ;
        RECT 164.910 125.600 165.750 125.880 ;
        RECT 153.990 125.320 157.070 125.600 ;
        RECT 122.070 124.480 125.150 124.760 ;
        RECT 125.990 125.040 128.790 125.320 ;
        RECT 131.590 125.040 131.870 125.320 ;
        RECT 135.230 125.040 137.470 125.320 ;
        RECT 140.550 125.040 141.670 125.320 ;
        RECT 142.790 125.040 143.630 125.320 ;
        RECT 146.990 125.040 147.270 125.320 ;
        RECT 151.470 125.040 152.870 125.320 ;
        RECT 125.990 124.480 128.510 125.040 ;
        RECT 131.590 124.760 132.150 125.040 ;
        RECT 135.510 124.760 137.190 125.040 ;
        RECT 140.830 124.760 141.670 125.040 ;
        RECT 142.510 124.760 143.350 125.040 ;
        RECT 146.710 124.760 147.270 125.040 ;
        RECT 122.070 123.640 125.430 124.480 ;
        RECT 126.270 123.640 128.230 124.480 ;
        RECT 131.870 124.200 132.430 124.760 ;
        RECT 135.790 124.480 136.910 124.760 ;
        RECT 140.830 124.480 143.070 124.760 ;
        RECT 146.710 124.480 146.990 124.760 ;
        RECT 136.070 124.200 137.190 124.480 ;
        RECT 141.110 124.200 142.790 124.480 ;
        RECT 146.430 124.200 146.990 124.480 ;
        RECT 151.190 124.200 152.870 125.040 ;
        RECT 153.710 124.480 157.070 125.320 ;
        RECT 161.550 125.040 162.670 125.600 ;
        RECT 164.630 125.320 165.750 125.600 ;
        RECT 166.030 125.600 167.150 125.880 ;
        RECT 164.630 125.040 165.470 125.320 ;
        RECT 161.270 124.480 162.390 125.040 ;
        RECT 164.350 124.480 165.470 125.040 ;
        RECT 166.030 124.760 166.870 125.600 ;
        RECT 167.430 125.320 168.270 125.880 ;
        RECT 168.830 125.600 171.630 125.880 ;
        RECT 171.770 125.740 178.630 125.880 ;
        RECT 171.910 125.600 178.630 125.740 ;
        RECT 168.550 125.320 169.950 125.600 ;
        RECT 170.090 125.460 171.350 125.600 ;
        RECT 170.230 125.320 171.350 125.460 ;
        RECT 171.910 125.320 174.430 125.600 ;
        RECT 167.150 125.040 169.670 125.320 ;
        RECT 170.230 125.040 171.070 125.320 ;
        RECT 171.630 125.040 174.430 125.320 ;
        RECT 174.710 125.320 176.390 125.600 ;
        RECT 176.950 125.320 178.070 125.600 ;
        RECT 190.110 125.320 193.470 125.880 ;
        RECT 194.310 125.600 202.990 126.160 ;
        RECT 204.110 125.600 204.670 126.160 ;
        RECT 207.190 125.600 208.030 126.160 ;
        RECT 208.590 125.880 210.550 126.160 ;
        RECT 208.870 125.600 210.270 125.880 ;
        RECT 211.110 125.600 211.950 126.160 ;
        RECT 219.230 125.880 220.070 126.160 ;
        RECT 221.470 125.880 222.590 126.160 ;
        RECT 219.790 125.600 220.350 125.880 ;
        RECT 222.030 125.600 223.150 125.880 ;
        RECT 194.030 125.320 203.270 125.600 ;
        RECT 204.390 125.320 204.950 125.600 ;
        RECT 174.710 125.040 176.110 125.320 ;
        RECT 176.950 125.040 177.510 125.320 ;
        RECT 167.150 124.760 169.390 125.040 ;
        RECT 169.950 124.760 171.070 125.040 ;
        RECT 171.910 124.760 174.150 125.040 ;
        RECT 189.830 124.760 193.190 125.320 ;
        RECT 193.750 125.040 203.270 125.320 ;
        RECT 204.670 125.040 204.950 125.320 ;
        RECT 207.470 125.320 208.310 125.600 ;
        RECT 210.830 125.320 211.670 125.600 ;
        RECT 220.070 125.320 220.910 125.600 ;
        RECT 222.310 125.320 223.430 125.600 ;
        RECT 207.470 125.040 208.870 125.320 ;
        RECT 210.270 125.040 211.390 125.320 ;
        RECT 220.350 125.040 221.190 125.320 ;
        RECT 222.590 125.040 223.710 125.320 ;
        RECT 193.750 124.760 203.550 125.040 ;
        RECT 204.670 124.760 205.230 125.040 ;
        RECT 207.750 124.760 211.110 125.040 ;
        RECT 220.910 124.760 221.750 125.040 ;
        RECT 222.870 124.760 223.990 125.040 ;
        RECT 165.750 124.480 167.710 124.760 ;
        RECT 167.990 124.480 169.110 124.760 ;
        RECT 170.230 124.480 170.790 124.760 ;
        RECT 172.610 124.620 173.870 124.760 ;
        RECT 172.750 124.480 173.870 124.620 ;
        RECT 189.550 124.480 192.910 124.760 ;
        RECT 193.470 124.480 203.550 124.760 ;
        RECT 204.950 124.480 205.230 124.760 ;
        RECT 208.310 124.480 210.830 124.760 ;
        RECT 221.190 124.480 222.030 124.760 ;
        RECT 223.430 124.480 224.270 124.760 ;
        RECT 132.150 123.920 132.710 124.200 ;
        RECT 136.630 123.920 138.030 124.200 ;
        RECT 140.830 123.920 142.510 124.200 ;
        RECT 122.350 123.080 125.710 123.640 ;
        RECT 126.550 123.080 128.230 123.640 ;
        RECT 132.430 123.360 132.990 123.920 ;
        RECT 136.910 123.640 141.950 123.920 ;
        RECT 146.150 123.640 146.710 124.200 ;
        RECT 150.910 123.640 152.590 124.200 ;
        RECT 153.430 123.640 156.790 124.480 ;
        RECT 160.990 124.200 162.110 124.480 ;
        RECT 160.710 123.920 161.830 124.200 ;
        RECT 137.750 123.360 141.390 123.640 ;
        RECT 145.870 123.360 146.430 123.640 ;
        RECT 132.710 123.080 133.270 123.360 ;
        RECT 145.590 123.080 146.430 123.360 ;
        RECT 150.630 123.080 152.310 123.640 ;
        RECT 122.350 122.800 125.990 123.080 ;
        RECT 122.630 122.520 125.990 122.800 ;
        RECT 126.830 122.800 128.510 123.080 ;
        RECT 132.990 122.800 133.550 123.080 ;
        RECT 145.310 122.800 146.710 123.080 ;
        RECT 126.830 122.520 128.790 122.800 ;
        RECT 133.270 122.520 133.830 122.800 ;
        RECT 145.030 122.520 146.710 122.800 ;
        RECT 150.350 122.800 152.310 123.080 ;
        RECT 153.150 123.360 156.790 123.640 ;
        RECT 160.430 123.640 161.830 123.920 ;
        RECT 164.070 123.920 165.190 124.480 ;
        RECT 165.750 123.920 167.430 124.480 ;
        RECT 168.270 124.200 168.550 124.480 ;
        RECT 172.470 124.200 173.870 124.480 ;
        RECT 172.190 123.920 173.590 124.200 ;
        RECT 178.630 123.920 178.910 124.200 ;
        RECT 189.270 123.920 192.630 124.480 ;
        RECT 193.470 124.200 203.830 124.480 ;
        RECT 204.950 124.200 205.510 124.480 ;
        RECT 209.150 124.200 209.990 124.480 ;
        RECT 221.750 124.200 222.310 124.480 ;
        RECT 223.710 124.200 224.550 124.480 ;
        RECT 193.190 123.920 204.110 124.200 ;
        RECT 164.070 123.640 164.910 123.920 ;
        RECT 165.750 123.640 167.150 123.920 ;
        RECT 171.910 123.640 173.030 123.920 ;
        RECT 178.070 123.640 178.350 123.920 ;
        RECT 188.990 123.640 192.350 123.920 ;
        RECT 192.910 123.640 204.110 123.920 ;
        RECT 205.230 123.920 205.510 124.200 ;
        RECT 222.030 123.920 222.870 124.200 ;
        RECT 223.990 123.920 225.110 124.200 ;
        RECT 205.230 123.640 205.790 123.920 ;
        RECT 222.310 123.640 223.150 123.920 ;
        RECT 224.270 123.640 225.390 123.920 ;
        RECT 240.510 123.640 241.350 123.920 ;
        RECT 160.430 123.360 162.110 123.640 ;
        RECT 164.070 123.360 164.630 123.640 ;
        RECT 165.750 123.360 166.870 123.640 ;
        RECT 171.630 123.360 172.190 123.640 ;
        RECT 177.510 123.360 177.790 123.640 ;
        RECT 153.150 122.800 156.510 123.360 ;
        RECT 160.430 123.080 162.950 123.360 ;
        RECT 171.350 123.080 171.910 123.360 ;
        RECT 176.670 123.080 177.230 123.360 ;
        RECT 188.710 123.080 192.070 123.640 ;
        RECT 192.910 123.360 204.390 123.640 ;
        RECT 205.510 123.360 205.790 123.640 ;
        RECT 222.870 123.360 223.710 123.640 ;
        RECT 224.550 123.360 225.670 123.640 ;
        RECT 192.630 123.080 200.470 123.360 ;
        RECT 202.430 123.080 204.670 123.360 ;
        RECT 205.510 123.080 206.070 123.360 ;
        RECT 223.150 123.080 223.990 123.360 ;
        RECT 225.110 123.080 225.950 123.360 ;
        RECT 240.230 123.080 241.630 123.640 ;
        RECT 160.990 122.800 163.790 123.080 ;
        RECT 170.790 122.940 171.490 123.080 ;
        RECT 175.830 122.940 176.810 123.080 ;
        RECT 170.790 122.800 171.350 122.940 ;
        RECT 175.830 122.800 176.670 122.940 ;
        RECT 188.430 122.800 191.790 123.080 ;
        RECT 192.350 122.800 199.910 123.080 ;
        RECT 200.750 122.800 204.670 123.080 ;
        RECT 205.790 122.800 206.070 123.080 ;
        RECT 223.710 122.800 224.270 123.080 ;
        RECT 225.390 122.800 226.230 123.080 ;
        RECT 150.350 122.520 152.030 122.800 ;
        RECT 122.630 121.960 126.270 122.520 ;
        RECT 127.110 122.240 128.790 122.520 ;
        RECT 133.550 122.240 134.110 122.520 ;
        RECT 144.750 122.240 146.990 122.520 ;
        RECT 150.070 122.240 152.030 122.520 ;
        RECT 152.870 122.520 156.510 122.800 ;
        RECT 161.830 122.520 164.630 122.800 ;
        RECT 170.790 122.520 171.070 122.800 ;
        RECT 174.710 122.660 175.970 122.800 ;
        RECT 174.710 122.520 175.830 122.660 ;
        RECT 152.870 122.240 156.230 122.520 ;
        RECT 162.670 122.240 165.750 122.520 ;
        RECT 173.590 122.240 174.990 122.520 ;
        RECT 188.150 122.240 191.510 122.800 ;
        RECT 192.350 122.520 199.630 122.800 ;
        RECT 200.190 122.520 201.030 122.800 ;
        RECT 202.150 122.520 204.950 122.800 ;
        RECT 205.930 122.660 206.350 122.800 ;
        RECT 127.110 121.960 129.070 122.240 ;
        RECT 133.830 121.960 134.670 122.240 ;
        RECT 144.190 121.960 145.030 122.240 ;
        RECT 145.590 121.960 146.990 122.240 ;
        RECT 149.790 121.960 151.750 122.240 ;
        RECT 152.590 121.960 156.230 122.240 ;
        RECT 163.510 121.960 167.710 122.240 ;
        RECT 171.630 121.960 173.870 122.240 ;
        RECT 187.870 121.960 191.230 122.240 ;
        RECT 192.070 121.960 199.350 122.520 ;
        RECT 199.910 122.240 200.470 122.520 ;
        RECT 202.710 122.240 205.230 122.520 ;
        RECT 206.070 122.240 206.350 122.660 ;
        RECT 223.990 122.520 224.830 122.800 ;
        RECT 225.670 122.520 226.510 122.800 ;
        RECT 239.950 122.520 241.910 123.080 ;
        RECT 224.270 122.240 225.110 122.520 ;
        RECT 225.950 122.240 226.790 122.520 ;
        RECT 199.910 121.960 200.190 122.240 ;
        RECT 122.910 121.400 126.550 121.960 ;
        RECT 127.390 121.680 129.070 121.960 ;
        RECT 134.390 121.680 134.950 121.960 ;
        RECT 143.910 121.680 144.750 121.960 ;
        RECT 145.590 121.680 147.550 121.960 ;
        RECT 149.510 121.680 151.470 121.960 ;
        RECT 152.590 121.680 155.950 121.960 ;
        RECT 164.910 121.680 172.750 121.960 ;
        RECT 187.590 121.680 191.230 121.960 ;
        RECT 191.790 121.680 199.070 121.960 ;
        RECT 127.390 121.400 129.350 121.680 ;
        RECT 134.670 121.400 135.510 121.680 ;
        RECT 143.350 121.400 144.190 121.680 ;
        RECT 145.590 121.400 148.110 121.680 ;
        RECT 148.950 121.400 151.470 121.680 ;
        RECT 152.310 121.400 155.950 121.680 ;
        RECT 167.150 121.400 170.510 121.680 ;
        RECT 187.590 121.400 190.950 121.680 ;
        RECT 123.190 120.840 126.830 121.400 ;
        RECT 127.670 121.120 129.630 121.400 ;
        RECT 135.230 121.120 136.070 121.400 ;
        RECT 142.790 121.120 143.910 121.400 ;
        RECT 145.590 121.120 151.190 121.400 ;
        RECT 123.470 120.560 127.110 120.840 ;
        RECT 127.950 120.560 129.910 121.120 ;
        RECT 135.790 120.840 136.910 121.120 ;
        RECT 142.230 120.840 143.350 121.120 ;
        RECT 145.870 120.840 151.190 121.120 ;
        RECT 152.030 121.120 155.950 121.400 ;
        RECT 152.030 120.840 155.670 121.120 ;
        RECT 187.310 120.840 190.670 121.400 ;
        RECT 191.510 121.120 199.070 121.680 ;
        RECT 191.230 120.840 199.070 121.120 ;
        RECT 136.350 120.560 137.750 120.840 ;
        RECT 141.110 120.560 142.510 120.840 ;
        RECT 145.870 120.560 150.910 120.840 ;
        RECT 151.750 120.560 155.670 120.840 ;
        RECT 187.030 120.560 190.390 120.840 ;
        RECT 191.230 120.560 193.750 120.840 ;
        RECT 123.470 120.280 127.390 120.560 ;
        RECT 128.230 120.280 130.190 120.560 ;
        RECT 137.190 120.280 141.670 120.560 ;
        RECT 145.870 120.280 150.630 120.560 ;
        RECT 151.750 120.280 155.390 120.560 ;
        RECT 123.750 120.000 127.390 120.280 ;
        RECT 128.510 120.000 130.470 120.280 ;
        RECT 138.590 120.000 140.550 120.280 ;
        RECT 123.750 119.720 127.670 120.000 ;
        RECT 128.790 119.720 130.750 120.000 ;
        RECT 138.870 119.720 140.550 120.000 ;
        RECT 145.870 119.720 150.350 120.280 ;
        RECT 151.470 120.000 155.110 120.280 ;
        RECT 186.750 120.000 190.110 120.560 ;
        RECT 191.790 120.280 193.470 120.560 ;
        RECT 192.350 120.000 193.470 120.280 ;
        RECT 151.190 119.720 155.110 120.000 ;
        RECT 186.470 119.720 189.830 120.000 ;
        RECT 192.910 119.720 193.190 120.000 ;
        RECT 195.150 119.720 199.070 120.840 ;
        RECT 199.630 121.680 200.190 121.960 ;
        RECT 202.990 121.960 205.510 122.240 ;
        RECT 224.550 121.960 225.390 122.240 ;
        RECT 226.230 121.960 227.070 122.240 ;
        RECT 239.670 121.960 242.190 122.520 ;
        RECT 202.990 121.820 203.690 121.960 ;
        RECT 202.990 121.680 203.550 121.820 ;
        RECT 199.630 120.840 199.910 121.680 ;
        RECT 203.270 120.840 203.550 121.680 ;
        RECT 199.630 120.560 200.190 120.840 ;
        RECT 199.910 120.280 200.190 120.560 ;
        RECT 202.990 120.560 203.550 120.840 ;
        RECT 203.830 121.400 205.790 121.960 ;
        RECT 225.110 121.680 225.950 121.960 ;
        RECT 226.510 121.680 227.350 121.960 ;
        RECT 239.670 121.680 242.470 121.960 ;
        RECT 225.390 121.400 226.230 121.680 ;
        RECT 226.790 121.400 227.630 121.680 ;
        RECT 239.670 121.400 242.750 121.680 ;
        RECT 203.830 121.120 206.070 121.400 ;
        RECT 225.670 121.120 226.510 121.400 ;
        RECT 227.070 121.120 227.910 121.400 ;
        RECT 239.670 121.120 243.030 121.400 ;
        RECT 203.830 120.840 206.350 121.120 ;
        RECT 225.950 120.840 226.790 121.120 ;
        RECT 227.350 120.840 228.470 121.120 ;
        RECT 203.830 120.560 206.630 120.840 ;
        RECT 226.510 120.560 228.750 120.840 ;
        RECT 239.670 120.560 242.470 121.120 ;
        RECT 242.750 120.840 243.030 121.120 ;
        RECT 242.750 120.560 243.310 120.840 ;
        RECT 202.990 120.280 203.270 120.560 ;
        RECT 199.910 120.000 200.470 120.280 ;
        RECT 202.710 120.000 203.270 120.280 ;
        RECT 203.830 120.280 206.910 120.560 ;
        RECT 226.790 120.420 227.770 120.560 ;
        RECT 226.790 120.280 227.630 120.420 ;
        RECT 228.190 120.280 229.030 120.560 ;
        RECT 203.830 120.000 207.190 120.280 ;
        RECT 227.070 120.000 227.910 120.280 ;
        RECT 228.470 120.000 229.030 120.280 ;
        RECT 239.670 120.420 242.890 120.560 ;
        RECT 200.190 119.720 200.750 120.000 ;
        RECT 202.430 119.720 202.990 120.000 ;
        RECT 203.550 119.720 207.470 120.000 ;
        RECT 227.350 119.720 228.190 120.000 ;
        RECT 239.670 119.720 242.750 120.420 ;
        RECT 243.030 120.280 243.310 120.560 ;
        RECT 243.030 120.000 243.590 120.280 ;
        RECT 124.030 119.440 127.950 119.720 ;
        RECT 129.070 119.440 131.030 119.720 ;
        RECT 124.310 119.160 128.230 119.440 ;
        RECT 129.070 119.160 131.590 119.440 ;
        RECT 138.870 119.160 140.830 119.720 ;
        RECT 124.310 118.880 128.510 119.160 ;
        RECT 129.350 118.880 131.870 119.160 ;
        RECT 139.150 118.880 140.830 119.160 ;
        RECT 146.150 119.440 150.070 119.720 ;
        RECT 150.910 119.440 154.830 119.720 ;
        RECT 146.150 119.160 149.790 119.440 ;
        RECT 150.630 119.160 154.830 119.440 ;
        RECT 186.190 119.440 189.830 119.720 ;
        RECT 186.190 119.160 189.550 119.440 ;
        RECT 146.150 118.880 149.510 119.160 ;
        RECT 150.630 118.880 154.550 119.160 ;
        RECT 185.910 118.880 189.270 119.160 ;
        RECT 124.590 118.600 128.790 118.880 ;
        RECT 129.630 118.600 132.150 118.880 ;
        RECT 124.870 118.320 128.790 118.600 ;
        RECT 129.910 118.320 132.710 118.600 ;
        RECT 139.150 118.320 141.110 118.880 ;
        RECT 146.150 118.600 149.230 118.880 ;
        RECT 150.350 118.600 154.270 118.880 ;
        RECT 146.150 118.320 148.950 118.600 ;
        RECT 150.070 118.320 154.270 118.600 ;
        RECT 185.630 118.600 189.270 118.880 ;
        RECT 195.430 118.600 198.790 119.720 ;
        RECT 200.470 119.440 202.710 119.720 ;
        RECT 203.550 119.440 208.030 119.720 ;
        RECT 227.630 119.440 228.470 119.720 ;
        RECT 238.270 119.440 242.750 119.720 ;
        RECT 201.310 119.160 201.870 119.440 ;
        RECT 203.550 119.160 208.310 119.440 ;
        RECT 228.190 119.160 229.030 119.440 ;
        RECT 237.710 119.160 242.750 119.440 ;
        RECT 185.630 118.320 188.990 118.600 ;
        RECT 124.870 118.040 129.350 118.320 ;
        RECT 130.470 118.040 132.990 118.320 ;
        RECT 139.150 118.040 141.390 118.320 ;
        RECT 145.870 118.040 148.670 118.320 ;
        RECT 149.790 118.040 153.990 118.320 ;
        RECT 185.350 118.040 188.710 118.320 ;
        RECT 125.150 117.760 129.630 118.040 ;
        RECT 130.750 117.760 133.550 118.040 ;
        RECT 138.870 117.760 141.390 118.040 ;
        RECT 145.310 117.760 148.110 118.040 ;
        RECT 149.510 117.760 153.710 118.040 ;
        RECT 185.070 117.760 188.710 118.040 ;
        RECT 195.710 118.040 198.790 118.600 ;
        RECT 203.550 118.880 209.150 119.160 ;
        RECT 228.470 118.880 229.310 119.160 ;
        RECT 237.430 118.880 239.670 119.160 ;
        RECT 239.950 118.880 242.750 119.160 ;
        RECT 243.310 119.720 243.590 120.000 ;
        RECT 243.310 118.880 243.870 119.720 ;
        RECT 203.550 118.600 210.550 118.880 ;
        RECT 228.750 118.600 229.590 118.880 ;
        RECT 237.150 118.600 238.830 118.880 ;
        RECT 203.550 118.320 207.750 118.600 ;
        RECT 208.590 118.320 211.950 118.600 ;
        RECT 229.030 118.320 229.870 118.600 ;
        RECT 202.990 118.040 207.750 118.320 ;
        RECT 209.430 118.040 213.630 118.320 ;
        RECT 229.310 118.040 230.150 118.320 ;
        RECT 237.150 118.040 238.270 118.600 ;
        RECT 240.230 118.320 242.750 118.880 ;
        RECT 239.950 118.040 242.750 118.320 ;
        RECT 125.430 117.480 129.910 117.760 ;
        RECT 131.030 117.480 134.110 117.760 ;
        RECT 125.710 117.200 130.190 117.480 ;
        RECT 131.310 117.200 134.670 117.480 ;
        RECT 138.870 117.200 141.670 117.760 ;
        RECT 144.750 117.480 147.830 117.760 ;
        RECT 148.950 117.480 153.430 117.760 ;
        RECT 185.070 117.480 188.430 117.760 ;
        RECT 194.590 117.480 194.870 117.760 ;
        RECT 144.190 117.200 147.550 117.480 ;
        RECT 148.670 117.200 153.430 117.480 ;
        RECT 184.790 117.200 188.430 117.480 ;
        RECT 193.750 117.200 195.150 117.480 ;
        RECT 195.710 117.200 198.510 118.040 ;
        RECT 202.430 117.760 207.750 118.040 ;
        RECT 211.110 117.760 215.030 118.040 ;
        RECT 229.590 117.760 230.150 118.040 ;
        RECT 201.870 117.480 206.350 117.760 ;
        RECT 212.790 117.480 216.710 117.760 ;
        RECT 237.430 117.480 238.270 118.040 ;
        RECT 201.030 117.200 204.950 117.480 ;
        RECT 213.350 117.200 218.390 117.480 ;
        RECT 237.710 117.200 238.270 117.480 ;
        RECT 238.830 117.760 239.390 118.040 ;
        RECT 240.510 117.760 242.750 118.040 ;
        RECT 243.590 118.600 243.870 118.880 ;
        RECT 125.710 116.920 130.470 117.200 ;
        RECT 131.870 116.920 135.510 117.200 ;
        RECT 138.590 116.920 141.950 117.200 ;
        RECT 143.350 116.920 146.990 117.200 ;
        RECT 148.390 116.920 153.150 117.200 ;
        RECT 184.790 116.920 188.150 117.200 ;
        RECT 192.630 117.060 193.890 117.200 ;
        RECT 192.630 116.920 193.750 117.060 ;
        RECT 194.590 116.920 195.430 117.200 ;
        RECT 195.990 116.920 198.230 117.200 ;
        RECT 199.910 116.920 203.270 117.200 ;
        RECT 209.150 116.920 211.670 117.200 ;
        RECT 213.630 116.920 214.750 117.200 ;
        RECT 216.150 116.920 219.790 117.200 ;
        RECT 125.990 116.640 131.030 116.920 ;
        RECT 132.430 116.640 136.350 116.920 ;
        RECT 138.030 116.640 141.950 116.920 ;
        RECT 142.510 116.640 146.710 116.920 ;
        RECT 148.110 116.640 152.870 116.920 ;
        RECT 184.510 116.640 187.870 116.920 ;
        RECT 191.790 116.640 192.910 116.920 ;
        RECT 194.870 116.640 201.870 116.920 ;
        RECT 207.750 116.640 211.950 116.920 ;
        RECT 126.270 116.360 131.310 116.640 ;
        RECT 132.710 116.360 146.150 116.640 ;
        RECT 147.550 116.360 152.590 116.640 ;
        RECT 184.230 116.360 187.870 116.640 ;
        RECT 190.950 116.500 191.930 116.640 ;
        RECT 190.950 116.360 191.790 116.500 ;
        RECT 194.870 116.360 200.470 116.640 ;
        RECT 206.630 116.360 212.230 116.640 ;
        RECT 213.910 116.360 215.030 116.920 ;
        RECT 217.830 116.640 221.470 116.920 ;
        RECT 237.710 116.640 238.550 117.200 ;
        RECT 238.830 116.920 239.110 117.760 ;
        RECT 240.790 117.480 242.470 117.760 ;
        RECT 241.070 117.200 242.470 117.480 ;
        RECT 238.970 116.780 239.390 116.920 ;
        RECT 219.510 116.360 222.870 116.640 ;
        RECT 126.550 116.080 131.870 116.360 ;
        RECT 133.270 116.080 145.590 116.360 ;
        RECT 147.270 116.080 152.310 116.360 ;
        RECT 184.230 116.080 187.590 116.360 ;
        RECT 190.670 116.220 191.090 116.360 ;
        RECT 126.830 115.800 132.150 116.080 ;
        RECT 134.110 115.800 145.030 116.080 ;
        RECT 146.710 115.800 152.030 116.080 ;
        RECT 183.950 115.800 187.310 116.080 ;
        RECT 127.110 115.520 132.710 115.800 ;
        RECT 134.670 115.520 144.190 115.800 ;
        RECT 146.150 115.520 151.750 115.800 ;
        RECT 183.670 115.520 187.310 115.800 ;
        RECT 127.390 115.240 133.270 115.520 ;
        RECT 135.510 115.240 143.350 115.520 ;
        RECT 145.590 115.240 151.470 115.520 ;
        RECT 183.670 115.240 187.030 115.520 ;
        RECT 190.670 115.240 190.950 116.220 ;
        RECT 194.870 115.800 199.910 116.360 ;
        RECT 205.790 116.080 209.990 116.360 ;
        RECT 211.110 116.080 212.230 116.360 ;
        RECT 204.670 115.800 209.150 116.080 ;
        RECT 193.190 115.520 194.590 115.800 ;
        RECT 192.350 115.380 193.330 115.520 ;
        RECT 192.350 115.240 193.190 115.380 ;
        RECT 127.950 114.960 134.110 115.240 ;
        RECT 136.630 114.960 142.230 115.240 ;
        RECT 145.030 114.960 151.190 115.240 ;
        RECT 167.150 114.960 173.590 115.240 ;
        RECT 183.390 114.960 187.030 115.240 ;
        RECT 190.810 115.100 191.230 115.240 ;
        RECT 128.230 114.680 134.670 114.960 ;
        RECT 144.190 114.680 150.630 114.960 ;
        RECT 165.750 114.680 174.990 114.960 ;
        RECT 183.110 114.680 186.750 114.960 ;
        RECT 128.510 114.400 135.790 114.680 ;
        RECT 143.350 114.400 150.350 114.680 ;
        RECT 164.630 114.400 167.430 114.680 ;
        RECT 173.310 114.400 176.110 114.680 ;
        RECT 183.110 114.400 186.470 114.680 ;
        RECT 128.790 114.120 136.910 114.400 ;
        RECT 141.950 114.120 150.070 114.400 ;
        RECT 164.070 114.120 166.030 114.400 ;
        RECT 174.710 114.120 177.230 114.400 ;
        RECT 182.830 114.120 186.470 114.400 ;
        RECT 190.950 114.120 191.230 115.100 ;
        RECT 192.350 114.400 192.630 115.240 ;
        RECT 194.310 114.680 194.590 115.520 ;
        RECT 195.150 115.520 199.910 115.800 ;
        RECT 203.830 115.520 209.150 115.800 ;
        RECT 211.110 115.800 212.510 116.080 ;
        RECT 214.190 115.800 215.310 116.360 ;
        RECT 221.190 116.080 224.550 116.360 ;
        RECT 222.870 115.800 225.950 116.080 ;
        RECT 237.990 115.800 238.830 116.640 ;
        RECT 239.110 116.080 239.390 116.780 ;
        RECT 241.350 116.640 242.190 117.200 ;
        RECT 241.630 116.360 242.470 116.640 ;
        RECT 243.590 116.360 244.150 118.600 ;
        RECT 241.910 116.080 242.750 116.360 ;
        RECT 243.310 116.080 244.150 116.360 ;
        RECT 239.250 115.940 239.670 116.080 ;
        RECT 195.150 115.240 200.190 115.520 ;
        RECT 202.990 115.240 208.870 115.520 ;
        RECT 211.110 115.240 212.790 115.800 ;
        RECT 214.190 115.520 215.590 115.800 ;
        RECT 224.550 115.520 227.070 115.800 ;
        RECT 214.470 115.240 215.590 115.520 ;
        RECT 225.950 115.240 227.630 115.520 ;
        RECT 238.270 115.240 239.110 115.800 ;
        RECT 239.390 115.240 239.670 115.940 ;
        RECT 241.910 115.800 243.870 116.080 ;
        RECT 242.190 115.520 243.870 115.800 ;
        RECT 242.750 115.240 243.590 115.520 ;
        RECT 195.150 114.960 201.590 115.240 ;
        RECT 195.150 114.680 201.870 114.960 ;
        RECT 202.710 114.680 208.590 115.240 ;
        RECT 211.390 114.960 213.070 115.240 ;
        RECT 211.110 114.680 213.070 114.960 ;
        RECT 214.470 114.680 215.870 115.240 ;
        RECT 227.070 114.960 227.630 115.240 ;
        RECT 238.550 115.100 239.950 115.240 ;
        RECT 194.450 114.540 194.870 114.680 ;
        RECT 192.490 114.260 192.910 114.400 ;
        RECT 129.350 113.840 149.510 114.120 ;
        RECT 163.510 113.840 165.190 114.120 ;
        RECT 175.830 113.840 178.070 114.120 ;
        RECT 182.550 113.840 186.190 114.120 ;
        RECT 191.090 113.980 191.510 114.120 ;
        RECT 129.630 113.560 149.230 113.840 ;
        RECT 163.230 113.560 164.350 113.840 ;
        RECT 176.670 113.560 178.630 113.840 ;
        RECT 182.550 113.560 185.910 113.840 ;
        RECT 130.190 113.280 148.670 113.560 ;
        RECT 163.230 113.280 164.070 113.560 ;
        RECT 177.510 113.280 179.470 113.560 ;
        RECT 182.270 113.280 185.910 113.560 ;
        RECT 130.750 113.000 148.390 113.280 ;
        RECT 163.510 113.000 164.630 113.280 ;
        RECT 178.350 113.000 180.030 113.280 ;
        RECT 182.270 113.000 185.630 113.280 ;
        RECT 191.230 113.000 191.510 113.980 ;
        RECT 192.630 113.280 192.910 114.260 ;
        RECT 194.590 113.560 194.870 114.540 ;
        RECT 195.430 113.560 201.870 114.680 ;
        RECT 202.430 114.400 204.110 114.680 ;
        RECT 205.510 114.400 208.310 114.680 ;
        RECT 210.550 114.400 213.350 114.680 ;
        RECT 202.430 114.120 203.550 114.400 ;
        RECT 206.070 114.120 208.310 114.400 ;
        RECT 209.430 114.120 213.350 114.400 ;
        RECT 202.430 113.840 203.270 114.120 ;
        RECT 194.730 113.420 195.150 113.560 ;
        RECT 192.770 113.140 193.190 113.280 ;
        RECT 131.030 112.720 147.830 113.000 ;
        RECT 163.790 112.720 165.750 113.000 ;
        RECT 179.190 112.720 180.590 113.000 ;
        RECT 181.990 112.720 185.630 113.000 ;
        RECT 191.370 112.860 191.790 113.000 ;
        RECT 131.590 112.440 147.270 112.720 ;
        RECT 164.070 112.440 167.430 112.720 ;
        RECT 179.750 112.440 181.150 112.720 ;
        RECT 181.710 112.440 185.350 112.720 ;
        RECT 132.430 112.160 146.710 112.440 ;
        RECT 163.230 112.160 169.670 112.440 ;
        RECT 180.310 112.160 185.070 112.440 ;
        RECT 132.990 111.880 145.870 112.160 ;
        RECT 162.390 111.880 171.630 112.160 ;
        RECT 180.870 111.880 185.070 112.160 ;
        RECT 191.510 111.880 191.790 112.860 ;
        RECT 192.910 112.160 193.190 113.140 ;
        RECT 194.870 112.440 195.150 113.420 ;
        RECT 195.710 112.720 202.150 113.560 ;
        RECT 202.430 113.280 203.550 113.840 ;
        RECT 206.630 113.560 213.630 114.120 ;
        RECT 214.750 113.560 216.150 114.680 ;
        RECT 238.550 114.400 239.390 115.100 ;
        RECT 239.670 114.400 239.950 115.100 ;
        RECT 238.830 114.260 240.230 114.400 ;
        RECT 238.830 113.840 239.670 114.260 ;
        RECT 239.110 113.560 239.670 113.840 ;
        RECT 239.950 113.560 240.230 114.260 ;
        RECT 206.350 113.280 213.910 113.560 ;
        RECT 202.430 113.000 203.830 113.280 ;
        RECT 205.510 113.000 208.310 113.280 ;
        RECT 195.010 112.300 195.430 112.440 ;
        RECT 193.050 112.020 193.470 112.160 ;
        RECT 133.830 111.600 145.030 111.880 ;
        RECT 161.830 111.600 173.030 111.880 ;
        RECT 181.150 111.600 184.790 111.880 ;
        RECT 191.650 111.740 192.070 111.880 ;
        RECT 134.670 111.320 144.190 111.600 ;
        RECT 161.270 111.320 174.150 111.600 ;
        RECT 181.150 111.320 184.510 111.600 ;
        RECT 136.070 111.040 143.070 111.320 ;
        RECT 160.710 111.040 174.990 111.320 ;
        RECT 180.870 111.040 184.510 111.320 ;
        RECT 191.790 111.040 192.070 111.740 ;
        RECT 193.190 111.040 193.470 112.020 ;
        RECT 195.150 111.320 195.430 112.300 ;
        RECT 195.990 112.160 202.150 112.720 ;
        RECT 202.710 112.720 203.830 113.000 ;
        RECT 204.670 112.720 206.910 113.000 ;
        RECT 195.990 111.600 202.430 112.160 ;
        RECT 202.710 111.600 207.190 112.720 ;
        RECT 207.750 112.160 208.310 113.000 ;
        RECT 208.870 113.000 213.910 113.280 ;
        RECT 208.870 112.720 212.790 113.000 ;
        RECT 213.350 112.720 213.910 113.000 ;
        RECT 214.750 112.720 216.430 113.560 ;
        RECT 218.390 112.720 223.150 113.000 ;
        RECT 234.910 112.720 238.550 113.560 ;
        RECT 239.110 113.000 240.510 113.560 ;
        RECT 239.390 112.720 240.510 113.000 ;
        RECT 260.950 112.720 261.790 115.240 ;
        RECT 263.750 114.400 264.590 115.240 ;
        RECT 263.470 113.560 264.310 114.400 ;
        RECT 265.710 114.120 266.550 115.240 ;
        RECT 267.670 114.120 269.070 115.240 ;
        RECT 270.750 114.400 271.590 115.240 ;
        RECT 273.830 114.960 275.790 115.240 ;
        RECT 277.470 114.960 280.270 115.240 ;
        RECT 273.550 114.680 276.070 114.960 ;
        RECT 265.430 113.840 266.550 114.120 ;
        RECT 263.190 112.720 264.030 113.560 ;
        RECT 265.430 112.720 266.270 113.840 ;
        RECT 267.390 113.560 269.070 114.120 ;
        RECT 267.390 112.720 268.230 113.560 ;
        RECT 208.870 112.440 211.670 112.720 ;
        RECT 212.650 112.580 214.190 112.720 ;
        RECT 212.790 112.440 214.190 112.580 ;
        RECT 214.750 112.440 224.830 112.720 ;
        RECT 209.150 112.160 210.550 112.440 ;
        RECT 211.530 112.300 213.350 112.440 ;
        RECT 211.670 112.160 213.350 112.300 ;
        RECT 214.750 112.160 218.950 112.440 ;
        RECT 222.870 112.160 225.670 112.440 ;
        RECT 207.750 111.880 208.590 112.160 ;
        RECT 209.150 111.880 209.430 112.160 ;
        RECT 210.410 112.020 211.950 112.160 ;
        RECT 210.550 111.880 211.950 112.020 ;
        RECT 214.190 111.880 216.990 112.160 ;
        RECT 224.550 111.880 225.390 112.160 ;
        RECT 208.030 111.600 208.310 111.880 ;
        RECT 209.290 111.740 210.830 111.880 ;
        RECT 209.430 111.600 210.830 111.740 ;
        RECT 214.470 111.600 215.590 111.880 ;
        RECT 195.290 111.180 195.710 111.320 ;
        RECT 138.030 110.760 140.830 111.040 ;
        RECT 160.150 110.760 176.110 111.040 ;
        RECT 159.590 110.480 176.670 110.760 ;
        RECT 180.590 110.480 184.230 111.040 ;
        RECT 191.790 110.760 192.350 111.040 ;
        RECT 193.330 110.900 193.750 111.040 ;
        RECT 159.030 110.200 177.510 110.480 ;
        RECT 180.310 110.200 184.510 110.480 ;
        RECT 158.750 109.920 178.070 110.200 ;
        RECT 180.030 109.920 184.790 110.200 ;
        RECT 192.070 109.920 192.350 110.760 ;
        RECT 193.470 109.920 193.750 110.900 ;
        RECT 195.430 110.200 195.710 111.180 ;
        RECT 196.270 110.480 202.430 111.600 ;
        RECT 202.990 111.320 207.190 111.600 ;
        RECT 208.170 111.460 209.710 111.600 ;
        RECT 208.310 111.320 209.710 111.460 ;
        RECT 212.790 111.320 214.190 111.600 ;
        RECT 202.990 111.040 206.070 111.320 ;
        RECT 207.050 111.180 208.590 111.320 ;
        RECT 207.190 111.040 208.590 111.180 ;
        RECT 211.670 111.040 214.190 111.320 ;
        RECT 214.470 111.320 215.030 111.600 ;
        RECT 202.990 110.760 204.950 111.040 ;
        RECT 205.930 110.900 207.470 111.040 ;
        RECT 206.070 110.760 207.470 110.900 ;
        RECT 210.550 110.760 213.070 111.040 ;
        RECT 214.470 110.760 215.310 111.320 ;
        RECT 202.990 110.480 203.830 110.760 ;
        RECT 204.810 110.620 206.350 110.760 ;
        RECT 204.950 110.480 206.350 110.620 ;
        RECT 209.430 110.480 211.950 110.760 ;
        RECT 213.350 110.620 214.610 110.760 ;
        RECT 213.350 110.480 214.470 110.620 ;
        RECT 195.570 110.060 195.990 110.200 ;
        RECT 158.190 109.640 178.630 109.920 ;
        RECT 180.030 109.640 183.670 109.920 ;
        RECT 184.230 109.640 185.070 109.920 ;
        RECT 192.210 109.780 192.630 109.920 ;
        RECT 193.610 109.780 194.030 109.920 ;
        RECT 157.910 109.360 167.150 109.640 ;
        RECT 172.750 109.360 179.190 109.640 ;
        RECT 179.750 109.360 183.390 109.640 ;
        RECT 184.510 109.360 185.350 109.640 ;
        RECT 157.630 109.080 165.750 109.360 ;
        RECT 174.150 109.080 183.110 109.360 ;
        RECT 184.790 109.080 185.630 109.360 ;
        RECT 157.070 108.800 164.910 109.080 ;
        RECT 174.990 108.800 183.110 109.080 ;
        RECT 185.070 108.800 185.910 109.080 ;
        RECT 192.350 108.800 192.630 109.780 ;
        RECT 193.750 108.800 194.030 109.780 ;
        RECT 195.710 109.080 195.990 110.060 ;
        RECT 196.550 109.360 202.710 110.480 ;
        RECT 203.270 110.200 205.230 110.480 ;
        RECT 208.310 110.200 210.830 110.480 ;
        RECT 212.230 110.200 214.470 110.480 ;
        RECT 214.750 110.200 215.310 110.760 ;
        RECT 234.910 110.480 235.190 112.720 ;
        RECT 236.870 112.160 237.430 112.440 ;
        RECT 236.590 111.880 237.710 112.160 ;
        RECT 237.990 111.880 238.270 112.720 ;
        RECT 239.390 112.440 240.790 112.720 ;
        RECT 236.590 111.600 236.870 111.880 ;
        RECT 237.570 111.740 238.270 111.880 ;
        RECT 237.710 111.600 238.270 111.740 ;
        RECT 239.670 111.880 240.790 112.440 ;
        RECT 239.670 111.600 241.070 111.880 ;
        RECT 236.310 111.460 236.730 111.600 ;
        RECT 236.310 111.320 236.590 111.460 ;
        RECT 237.990 111.320 238.550 111.600 ;
        RECT 236.030 111.040 236.590 111.320 ;
        RECT 238.270 111.040 239.110 111.320 ;
        RECT 239.950 111.040 241.070 111.600 ;
        RECT 242.750 111.320 244.710 111.600 ;
        RECT 242.190 111.040 245.270 111.320 ;
        RECT 245.830 111.040 247.230 111.320 ;
        RECT 235.750 110.760 236.310 111.040 ;
        RECT 237.710 110.900 238.410 111.040 ;
        RECT 237.710 110.760 238.270 110.900 ;
        RECT 238.830 110.760 239.390 111.040 ;
        RECT 240.230 110.760 241.350 111.040 ;
        RECT 241.910 110.760 247.790 111.040 ;
        RECT 235.750 110.480 236.030 110.760 ;
        RECT 237.430 110.480 237.990 110.760 ;
        RECT 239.250 110.620 239.950 110.760 ;
        RECT 239.390 110.480 239.950 110.620 ;
        RECT 240.230 110.480 246.110 110.760 ;
        RECT 247.230 110.480 248.070 110.760 ;
        RECT 235.050 110.340 235.890 110.480 ;
        RECT 235.190 110.200 235.750 110.340 ;
        RECT 237.430 110.200 237.710 110.480 ;
        RECT 239.670 110.200 245.550 110.480 ;
        RECT 203.270 109.920 204.110 110.200 ;
        RECT 207.190 109.920 209.990 110.200 ;
        RECT 211.110 109.920 213.910 110.200 ;
        RECT 206.070 109.640 208.870 109.920 ;
        RECT 210.270 109.640 212.790 109.920 ;
        RECT 214.190 109.640 214.470 109.920 ;
        RECT 214.750 109.640 215.590 110.200 ;
        RECT 235.190 109.920 235.470 110.200 ;
        RECT 237.150 110.060 237.570 110.200 ;
        RECT 237.150 109.920 237.430 110.060 ;
        RECT 240.230 109.920 244.990 110.200 ;
        RECT 225.670 109.640 226.790 109.920 ;
        RECT 234.910 109.640 235.470 109.920 ;
        RECT 236.870 109.780 237.290 109.920 ;
        RECT 236.870 109.640 237.150 109.780 ;
        RECT 240.510 109.640 244.430 109.920 ;
        RECT 204.950 109.360 207.750 109.640 ;
        RECT 209.150 109.360 211.670 109.640 ;
        RECT 213.070 109.500 214.890 109.640 ;
        RECT 213.070 109.360 214.750 109.500 ;
        RECT 196.830 109.080 201.870 109.360 ;
        RECT 204.110 109.080 206.630 109.360 ;
        RECT 208.030 109.080 210.550 109.360 ;
        RECT 211.950 109.080 214.470 109.360 ;
        RECT 215.030 109.080 215.590 109.640 ;
        RECT 225.390 109.360 227.070 109.640 ;
        RECT 234.910 109.360 235.190 109.640 ;
        RECT 236.590 109.360 237.150 109.640 ;
        RECT 240.790 109.360 243.870 109.640 ;
        RECT 247.510 109.360 248.070 110.480 ;
        RECT 260.670 109.640 261.510 112.720 ;
        RECT 262.910 111.880 263.750 112.720 ;
        RECT 262.630 111.320 263.470 111.880 ;
        RECT 265.150 111.320 265.990 112.720 ;
        RECT 267.110 111.320 267.950 112.720 ;
        RECT 262.630 111.040 263.190 111.320 ;
        RECT 262.350 110.480 263.190 111.040 ;
        RECT 262.070 109.640 262.910 110.480 ;
        RECT 264.870 110.200 265.710 111.320 ;
        RECT 266.830 110.200 267.670 111.320 ;
        RECT 264.590 109.920 265.710 110.200 ;
        RECT 266.550 109.920 267.670 110.200 ;
        RECT 216.990 109.080 221.470 109.360 ;
        RECT 225.110 109.080 225.950 109.360 ;
        RECT 226.510 109.080 227.350 109.360 ;
        RECT 234.630 109.220 235.050 109.360 ;
        RECT 234.630 109.080 234.910 109.220 ;
        RECT 236.590 109.080 236.870 109.360 ;
        RECT 238.550 109.080 242.470 109.360 ;
        RECT 247.230 109.080 247.790 109.360 ;
        RECT 260.670 109.080 261.230 109.640 ;
        RECT 195.850 108.940 196.270 109.080 ;
        RECT 156.790 108.520 164.070 108.800 ;
        RECT 167.710 108.520 172.190 108.800 ;
        RECT 175.830 108.520 182.830 108.800 ;
        RECT 185.350 108.520 186.190 108.800 ;
        RECT 192.490 108.660 192.910 108.800 ;
        RECT 193.890 108.660 194.310 108.800 ;
        RECT 156.510 108.240 163.230 108.520 ;
        RECT 166.030 108.240 173.870 108.520 ;
        RECT 176.670 108.240 182.550 108.520 ;
        RECT 185.630 108.240 186.470 108.520 ;
        RECT 156.230 107.960 162.670 108.240 ;
        RECT 165.190 107.960 174.710 108.240 ;
        RECT 177.230 107.960 182.550 108.240 ;
        RECT 185.910 107.960 186.750 108.240 ;
        RECT 155.950 107.680 162.110 107.960 ;
        RECT 164.350 107.680 175.550 107.960 ;
        RECT 177.790 107.680 182.270 107.960 ;
        RECT 186.190 107.680 187.030 107.960 ;
        RECT 192.630 107.680 192.910 108.660 ;
        RECT 194.030 107.680 194.310 108.660 ;
        RECT 195.990 107.960 196.270 108.940 ;
        RECT 196.830 108.240 200.750 109.080 ;
        RECT 196.130 107.820 196.550 107.960 ;
        RECT 155.670 107.400 161.550 107.680 ;
        RECT 163.510 107.400 176.390 107.680 ;
        RECT 178.350 107.400 182.550 107.680 ;
        RECT 186.470 107.400 187.030 107.680 ;
        RECT 192.770 107.540 193.190 107.680 ;
        RECT 194.170 107.540 194.590 107.680 ;
        RECT 155.390 107.120 161.270 107.400 ;
        RECT 162.950 107.120 176.950 107.400 ;
        RECT 178.350 107.120 182.830 107.400 ;
        RECT 186.470 107.120 187.310 107.400 ;
        RECT 155.110 106.840 160.710 107.120 ;
        RECT 162.390 106.840 177.510 107.120 ;
        RECT 178.070 106.840 183.110 107.120 ;
        RECT 186.750 106.840 187.590 107.120 ;
        RECT 154.830 106.560 160.430 106.840 ;
        RECT 161.830 106.560 166.590 106.840 ;
        RECT 167.710 106.560 171.910 106.840 ;
        RECT 173.310 106.560 183.390 106.840 ;
        RECT 154.550 106.280 159.870 106.560 ;
        RECT 161.550 106.280 165.750 106.560 ;
        RECT 154.270 106.000 159.590 106.280 ;
        RECT 160.990 106.000 164.910 106.280 ;
        RECT 167.990 106.000 169.670 106.560 ;
        RECT 153.990 105.720 159.310 106.000 ;
        RECT 160.710 105.720 164.350 106.000 ;
        RECT 168.270 105.720 169.670 106.000 ;
        RECT 153.710 105.440 158.750 105.720 ;
        RECT 160.150 105.440 163.510 105.720 ;
        RECT 153.710 105.160 158.470 105.440 ;
        RECT 159.870 105.160 163.230 105.440 ;
        RECT 168.550 105.160 169.670 105.720 ;
        RECT 153.430 104.880 158.190 105.160 ;
        RECT 159.590 104.880 162.670 105.160 ;
        RECT 153.150 104.600 157.910 104.880 ;
        RECT 159.310 104.600 162.110 104.880 ;
        RECT 152.870 104.320 157.630 104.600 ;
        RECT 159.030 104.320 161.830 104.600 ;
        RECT 152.870 104.040 157.350 104.320 ;
        RECT 158.750 104.040 161.270 104.320 ;
        RECT 152.590 103.760 157.070 104.040 ;
        RECT 158.470 103.760 160.990 104.040 ;
        RECT 152.310 103.480 157.070 103.760 ;
        RECT 158.190 103.480 160.710 103.760 ;
        RECT 152.310 103.200 156.790 103.480 ;
        RECT 157.910 103.200 160.430 103.480 ;
        RECT 168.830 103.200 169.670 105.160 ;
        RECT 152.030 102.920 156.510 103.200 ;
        RECT 157.630 102.920 160.150 103.200 ;
        RECT 152.030 102.640 156.230 102.920 ;
        RECT 157.350 102.640 159.870 102.920 ;
        RECT 151.750 102.360 156.230 102.640 ;
        RECT 157.070 102.360 159.590 102.640 ;
        RECT 151.750 102.080 155.950 102.360 ;
        RECT 157.070 102.080 159.310 102.360 ;
        RECT 169.110 102.080 169.670 103.200 ;
        RECT 169.950 106.280 171.630 106.560 ;
        RECT 174.150 106.280 183.670 106.560 ;
        RECT 187.030 106.280 187.870 106.840 ;
        RECT 192.910 106.560 193.190 107.540 ;
        RECT 194.310 106.840 194.590 107.540 ;
        RECT 196.270 106.840 196.550 107.820 ;
        RECT 197.110 107.400 200.750 108.240 ;
        RECT 201.590 108.800 201.870 109.080 ;
        RECT 202.990 108.800 205.510 109.080 ;
        RECT 206.910 108.800 209.430 109.080 ;
        RECT 210.830 108.800 213.350 109.080 ;
        RECT 215.030 108.800 221.470 109.080 ;
        RECT 224.830 108.800 225.670 109.080 ;
        RECT 226.790 108.800 227.630 109.080 ;
        RECT 234.350 108.940 234.770 109.080 ;
        RECT 234.350 108.800 234.630 108.940 ;
        RECT 235.750 108.800 240.510 109.080 ;
        RECT 246.950 108.800 247.790 109.080 ;
        RECT 201.590 108.520 204.390 108.800 ;
        RECT 205.790 108.520 208.310 108.800 ;
        RECT 209.710 108.520 212.230 108.800 ;
        RECT 213.630 108.520 214.750 108.800 ;
        RECT 215.030 108.520 217.550 108.800 ;
        RECT 220.910 108.520 221.190 108.800 ;
        RECT 201.590 108.240 203.270 108.520 ;
        RECT 204.670 108.240 207.190 108.520 ;
        RECT 208.590 108.240 211.110 108.520 ;
        RECT 212.510 108.240 214.750 108.520 ;
        RECT 215.310 108.240 215.870 108.520 ;
        RECT 224.830 108.240 225.390 108.800 ;
        RECT 227.070 108.520 227.910 108.800 ;
        RECT 234.070 108.520 238.270 108.800 ;
        RECT 246.390 108.520 247.510 108.800 ;
        RECT 227.350 108.240 228.190 108.520 ;
        RECT 233.790 108.240 235.470 108.520 ;
        RECT 245.830 108.240 247.230 108.520 ;
        RECT 201.590 107.960 202.150 108.240 ;
        RECT 203.550 107.960 206.070 108.240 ;
        RECT 207.470 107.960 209.990 108.240 ;
        RECT 211.390 107.960 213.910 108.240 ;
        RECT 216.430 107.960 216.990 108.240 ;
        RECT 224.830 107.960 225.670 108.240 ;
        RECT 227.630 107.960 228.470 108.240 ;
        RECT 233.230 107.960 234.630 108.240 ;
        RECT 244.990 107.960 246.670 108.240 ;
        RECT 201.870 107.680 202.150 107.960 ;
        RECT 202.430 107.680 204.950 107.960 ;
        RECT 206.350 107.680 208.870 107.960 ;
        RECT 210.270 107.680 212.790 107.960 ;
        RECT 215.310 107.680 218.110 107.960 ;
        RECT 225.110 107.680 225.670 107.960 ;
        RECT 227.910 107.680 228.750 107.960 ;
        RECT 233.230 107.680 234.070 107.960 ;
        RECT 243.870 107.680 246.110 107.960 ;
        RECT 201.870 107.400 203.830 107.680 ;
        RECT 205.230 107.400 207.750 107.680 ;
        RECT 209.150 107.400 211.670 107.680 ;
        RECT 214.750 107.400 215.590 107.680 ;
        RECT 217.830 107.400 218.390 107.680 ;
        RECT 225.110 107.400 225.950 107.680 ;
        RECT 228.190 107.400 229.030 107.680 ;
        RECT 197.390 107.120 200.470 107.400 ;
        RECT 201.870 107.120 202.710 107.400 ;
        RECT 204.110 107.120 206.630 107.400 ;
        RECT 208.030 107.120 210.550 107.400 ;
        RECT 214.470 107.120 215.030 107.400 ;
        RECT 218.110 107.120 218.670 107.400 ;
        RECT 224.830 107.120 226.230 107.400 ;
        RECT 228.470 107.120 229.030 107.400 ;
        RECT 197.390 106.840 200.190 107.120 ;
        RECT 201.310 106.840 202.150 107.120 ;
        RECT 202.990 106.840 205.510 107.120 ;
        RECT 206.910 106.840 209.710 107.120 ;
        RECT 214.190 106.840 214.750 107.120 ;
        RECT 218.530 106.980 218.950 107.120 ;
        RECT 218.670 106.840 218.950 106.980 ;
        RECT 194.310 106.560 194.870 106.840 ;
        RECT 196.410 106.700 196.830 106.840 ;
        RECT 193.050 106.420 193.470 106.560 ;
        RECT 169.950 106.000 171.350 106.280 ;
        RECT 174.990 106.000 183.950 106.280 ;
        RECT 187.310 106.000 188.150 106.280 ;
        RECT 169.950 105.440 171.070 106.000 ;
        RECT 175.550 105.720 184.230 106.000 ;
        RECT 187.590 105.720 188.150 106.000 ;
        RECT 176.390 105.440 184.510 105.720 ;
        RECT 187.590 105.440 188.430 105.720 ;
        RECT 193.190 105.440 193.470 106.420 ;
        RECT 194.590 105.720 194.870 106.560 ;
        RECT 196.550 106.000 196.830 106.700 ;
        RECT 197.390 106.560 199.910 106.840 ;
        RECT 200.750 106.560 201.870 106.840 ;
        RECT 202.010 106.700 204.670 106.840 ;
        RECT 197.390 106.280 199.350 106.560 ;
        RECT 200.470 106.280 201.870 106.560 ;
        RECT 195.710 105.720 196.830 106.000 ;
        RECT 197.670 106.000 199.070 106.280 ;
        RECT 199.910 106.000 200.750 106.280 ;
        RECT 201.310 106.000 201.870 106.280 ;
        RECT 197.670 105.720 198.790 106.000 ;
        RECT 199.630 105.720 200.470 106.000 ;
        RECT 201.590 105.720 201.870 106.000 ;
        RECT 202.150 106.560 204.670 106.700 ;
        RECT 205.790 106.560 208.590 106.840 ;
        RECT 213.910 106.560 214.470 106.840 ;
        RECT 218.670 106.560 219.230 106.840 ;
        RECT 224.830 106.560 225.390 107.120 ;
        RECT 225.670 106.840 226.510 107.120 ;
        RECT 228.750 106.840 229.310 107.120 ;
        RECT 233.230 106.840 233.790 107.680 ;
        RECT 242.190 107.400 246.110 107.680 ;
        RECT 239.110 107.120 246.110 107.400 ;
        RECT 236.030 106.840 246.110 107.120 ;
        RECT 260.390 107.680 261.230 109.080 ;
        RECT 261.790 108.800 262.630 109.640 ;
        RECT 264.590 108.800 265.430 109.920 ;
        RECT 266.550 108.800 267.390 109.920 ;
        RECT 261.510 107.960 262.350 108.800 ;
        RECT 261.510 107.680 262.070 107.960 ;
        RECT 260.390 107.120 262.070 107.680 ;
        RECT 264.310 107.400 265.150 108.800 ;
        RECT 266.270 107.400 267.110 108.800 ;
        RECT 268.510 108.520 269.070 113.560 ;
        RECT 270.470 114.120 271.590 114.400 ;
        RECT 272.990 114.400 276.070 114.680 ;
        RECT 277.470 114.400 279.990 114.960 ;
        RECT 272.990 114.120 274.110 114.400 ;
        RECT 270.470 113.000 271.310 114.120 ;
        RECT 272.710 113.840 273.830 114.120 ;
        RECT 272.710 113.000 273.550 113.840 ;
        RECT 270.190 112.720 271.310 113.000 ;
        RECT 272.430 112.720 273.550 113.000 ;
        RECT 275.230 113.560 276.350 114.400 ;
        RECT 277.470 114.120 278.310 114.400 ;
        RECT 281.390 114.120 282.790 115.240 ;
        RECT 284.470 114.400 285.310 115.240 ;
        RECT 286.150 114.960 289.230 115.240 ;
        RECT 291.750 114.960 294.550 115.240 ;
        RECT 285.870 114.400 288.950 114.960 ;
        RECT 291.750 114.400 294.270 114.960 ;
        RECT 277.190 113.840 278.310 114.120 ;
        RECT 270.190 111.600 271.030 112.720 ;
        RECT 272.430 111.600 273.270 112.720 ;
        RECT 275.230 112.440 276.070 113.560 ;
        RECT 277.190 112.720 278.030 113.840 ;
        RECT 281.110 113.560 282.790 114.120 ;
        RECT 281.110 112.720 281.950 113.560 ;
        RECT 274.950 112.160 275.790 112.440 ;
        RECT 276.910 111.600 277.750 112.720 ;
        RECT 269.910 110.480 270.750 111.600 ;
        RECT 269.630 110.200 270.750 110.480 ;
        RECT 272.150 110.200 272.990 111.600 ;
        RECT 276.910 111.320 279.150 111.600 ;
        RECT 280.830 111.320 281.670 112.720 ;
        RECT 276.630 110.760 279.150 111.320 ;
        RECT 276.630 110.200 277.470 110.760 ;
        RECT 280.550 110.200 281.390 111.320 ;
        RECT 269.630 108.800 270.470 110.200 ;
        RECT 271.870 109.080 272.710 110.200 ;
        RECT 276.350 109.920 277.470 110.200 ;
        RECT 280.270 109.920 281.390 110.200 ;
        RECT 271.590 108.800 272.710 109.080 ;
        RECT 274.390 109.640 275.510 109.920 ;
        RECT 269.350 108.520 270.190 108.800 ;
        RECT 268.510 107.680 270.190 108.520 ;
        RECT 271.590 107.960 272.430 108.800 ;
        RECT 274.390 108.520 275.230 109.640 ;
        RECT 276.350 108.800 277.190 109.920 ;
        RECT 280.270 108.800 281.110 109.920 ;
        RECT 274.110 108.240 275.230 108.520 ;
        RECT 274.110 107.960 274.950 108.240 ;
        RECT 271.590 107.680 272.710 107.960 ;
        RECT 273.830 107.680 274.950 107.960 ;
        RECT 276.070 107.680 276.910 108.800 ;
        RECT 260.390 106.840 261.790 107.120 ;
        RECT 264.030 106.840 264.870 107.400 ;
        RECT 265.990 106.840 266.830 107.400 ;
        RECT 268.510 106.840 269.910 107.680 ;
        RECT 271.590 107.400 274.670 107.680 ;
        RECT 276.070 107.400 278.590 107.680 ;
        RECT 279.990 107.400 280.830 108.800 ;
        RECT 282.230 108.520 282.790 113.560 ;
        RECT 284.190 114.120 285.310 114.400 ;
        RECT 284.190 113.000 285.030 114.120 ;
        RECT 286.990 113.560 287.830 114.400 ;
        RECT 291.750 114.120 292.590 114.400 ;
        RECT 295.390 114.120 296.230 115.240 ;
        RECT 298.190 114.960 299.030 115.240 ;
        RECT 300.710 114.960 302.670 115.240 ;
        RECT 305.470 114.960 307.430 115.240 ;
        RECT 309.950 114.960 311.910 115.240 ;
        RECT 291.470 113.840 292.590 114.120 ;
        RECT 283.910 112.720 285.030 113.000 ;
        RECT 283.910 111.600 284.750 112.720 ;
        RECT 286.710 112.440 287.550 113.560 ;
        RECT 291.470 112.720 292.310 113.840 ;
        RECT 295.110 112.720 295.950 114.120 ;
        RECT 297.910 113.560 298.750 114.960 ;
        RECT 300.430 114.680 302.950 114.960 ;
        RECT 305.190 114.680 307.710 114.960 ;
        RECT 309.670 114.680 312.190 114.960 ;
        RECT 300.150 114.400 303.230 114.680 ;
        RECT 299.870 114.120 300.990 114.400 ;
        RECT 302.110 114.120 303.230 114.400 ;
        RECT 304.630 114.400 307.710 114.680 ;
        RECT 309.110 114.400 312.190 114.680 ;
        RECT 304.630 114.120 305.750 114.400 ;
        RECT 299.870 113.560 300.710 114.120 ;
        RECT 286.430 112.160 287.550 112.440 ;
        RECT 283.630 110.480 284.470 111.600 ;
        RECT 286.430 111.040 287.270 112.160 ;
        RECT 291.190 111.600 292.030 112.720 ;
        RECT 294.830 111.600 295.670 112.720 ;
        RECT 297.630 112.440 298.470 113.560 ;
        RECT 299.590 112.440 300.430 113.560 ;
        RECT 302.390 113.280 303.230 114.120 ;
        RECT 304.350 113.840 305.470 114.120 ;
        RECT 302.110 112.720 302.950 113.280 ;
        RECT 304.350 113.000 305.190 113.840 ;
        RECT 304.070 112.720 305.190 113.000 ;
        RECT 306.870 113.560 307.990 114.400 ;
        RECT 309.110 114.120 310.230 114.400 ;
        RECT 308.830 113.840 309.950 114.120 ;
        RECT 291.190 111.320 293.430 111.600 ;
        RECT 283.350 110.200 284.470 110.480 ;
        RECT 286.150 110.760 287.270 111.040 ;
        RECT 290.910 110.760 293.430 111.320 ;
        RECT 294.550 111.320 295.670 111.600 ;
        RECT 297.350 112.160 298.470 112.440 ;
        RECT 299.310 112.160 300.430 112.440 ;
        RECT 283.350 108.800 284.190 110.200 ;
        RECT 286.150 109.640 286.990 110.760 ;
        RECT 290.910 110.200 291.750 110.760 ;
        RECT 294.550 110.200 295.390 111.320 ;
        RECT 297.350 111.040 298.190 112.160 ;
        RECT 299.310 111.880 300.710 112.160 ;
        RECT 299.590 111.600 300.990 111.880 ;
        RECT 304.070 111.600 304.910 112.720 ;
        RECT 306.870 112.440 307.710 113.560 ;
        RECT 308.830 113.000 309.670 113.840 ;
        RECT 308.550 112.720 309.670 113.000 ;
        RECT 311.350 113.560 312.470 114.400 ;
        RECT 306.590 112.160 307.430 112.440 ;
        RECT 308.550 111.600 309.390 112.720 ;
        RECT 311.350 112.440 312.190 113.560 ;
        RECT 299.870 111.320 301.270 111.600 ;
        RECT 300.150 111.040 301.550 111.320 ;
        RECT 290.630 109.920 291.750 110.200 ;
        RECT 283.070 108.520 283.910 108.800 ;
        RECT 282.230 107.680 283.910 108.520 ;
        RECT 285.870 108.240 286.710 109.640 ;
        RECT 290.630 108.800 291.470 109.920 ;
        RECT 294.270 108.800 295.110 110.200 ;
        RECT 297.070 109.640 297.910 111.040 ;
        RECT 300.430 110.760 301.830 111.040 ;
        RECT 300.710 110.480 302.110 110.760 ;
        RECT 300.990 110.200 302.390 110.480 ;
        RECT 303.790 110.200 304.630 111.600 ;
        RECT 308.270 110.200 309.110 111.600 ;
        RECT 311.070 111.040 311.910 112.440 ;
        RECT 301.270 109.920 302.390 110.200 ;
        RECT 271.870 107.120 274.390 107.400 ;
        RECT 272.150 106.840 274.110 107.120 ;
        RECT 275.790 106.840 278.590 107.400 ;
        RECT 279.710 106.840 280.550 107.400 ;
        RECT 282.230 106.840 283.630 107.680 ;
        RECT 285.590 107.120 286.430 108.240 ;
        RECT 290.350 107.400 291.190 108.800 ;
        RECT 293.990 107.960 294.830 108.800 ;
        RECT 296.790 108.520 297.630 109.640 ;
        RECT 298.750 108.520 299.590 109.640 ;
        RECT 301.550 109.360 302.390 109.920 ;
        RECT 296.510 108.240 297.630 108.520 ;
        RECT 296.510 107.960 297.350 108.240 ;
        RECT 293.990 107.680 295.110 107.960 ;
        RECT 296.230 107.680 297.350 107.960 ;
        RECT 298.470 107.680 299.590 108.520 ;
        RECT 301.270 109.080 302.390 109.360 ;
        RECT 303.510 109.080 304.350 110.200 ;
        RECT 301.270 108.240 302.110 109.080 ;
        RECT 300.990 107.960 302.110 108.240 ;
        RECT 303.230 108.800 304.350 109.080 ;
        RECT 306.030 109.640 307.150 109.920 ;
        RECT 303.230 107.960 304.070 108.800 ;
        RECT 306.030 108.520 306.870 109.640 ;
        RECT 307.990 109.080 308.830 110.200 ;
        RECT 310.790 109.920 311.630 111.040 ;
        RECT 305.750 108.240 306.870 108.520 ;
        RECT 307.710 108.800 308.830 109.080 ;
        RECT 310.510 109.640 311.630 109.920 ;
        RECT 305.750 107.960 306.590 108.240 ;
        RECT 300.710 107.680 301.830 107.960 ;
        RECT 293.990 107.400 297.070 107.680 ;
        RECT 298.750 107.400 301.830 107.680 ;
        RECT 303.230 107.680 304.350 107.960 ;
        RECT 305.470 107.680 306.590 107.960 ;
        RECT 307.710 107.960 308.550 108.800 ;
        RECT 310.510 108.520 311.350 109.640 ;
        RECT 310.230 108.240 311.350 108.520 ;
        RECT 310.230 107.960 311.070 108.240 ;
        RECT 307.710 107.680 308.830 107.960 ;
        RECT 309.950 107.680 311.070 107.960 ;
        RECT 303.230 107.400 306.310 107.680 ;
        RECT 307.710 107.400 310.790 107.680 ;
        RECT 285.310 106.840 286.430 107.120 ;
        RECT 290.070 106.840 290.910 107.400 ;
        RECT 294.270 107.120 296.790 107.400 ;
        RECT 298.750 107.120 301.270 107.400 ;
        RECT 303.510 107.120 306.030 107.400 ;
        RECT 307.990 107.120 310.510 107.400 ;
        RECT 294.550 106.840 296.510 107.120 ;
        RECT 299.030 106.840 300.990 107.120 ;
        RECT 303.790 106.840 305.750 107.120 ;
        RECT 308.270 106.840 310.230 107.120 ;
        RECT 225.950 106.560 226.790 106.840 ;
        RECT 228.750 106.560 229.590 106.840 ;
        RECT 202.150 106.280 203.550 106.560 ;
        RECT 204.530 106.420 207.470 106.560 ;
        RECT 204.670 106.280 207.470 106.420 ;
        RECT 209.150 106.280 209.990 106.560 ;
        RECT 210.830 106.280 211.390 106.560 ;
        RECT 213.910 106.280 214.190 106.560 ;
        RECT 218.950 106.280 219.510 106.560 ;
        RECT 224.830 106.280 225.670 106.560 ;
        RECT 225.950 106.280 227.070 106.560 ;
        RECT 229.030 106.280 229.870 106.560 ;
        RECT 233.510 106.280 234.070 106.840 ;
        RECT 235.750 106.560 238.270 106.840 ;
        RECT 241.630 106.560 246.110 106.840 ;
        RECT 235.470 106.280 236.310 106.560 ;
        RECT 241.350 106.280 246.110 106.560 ;
        RECT 202.150 106.000 202.430 106.280 ;
        RECT 203.830 106.000 206.350 106.280 ;
        RECT 208.030 106.000 208.870 106.280 ;
        RECT 211.250 106.140 212.230 106.280 ;
        RECT 211.390 106.000 212.230 106.140 ;
        RECT 202.150 105.720 205.230 106.000 ;
        RECT 207.190 105.720 207.750 106.000 ;
        RECT 210.550 105.720 212.230 106.000 ;
        RECT 213.630 106.000 214.190 106.280 ;
        RECT 194.730 105.580 195.850 105.720 ;
        RECT 194.870 105.440 195.710 105.580 ;
        RECT 197.670 105.440 198.510 105.720 ;
        RECT 199.350 105.440 200.190 105.720 ;
        RECT 201.590 105.580 202.290 105.720 ;
        RECT 169.950 104.880 170.790 105.440 ;
        RECT 176.670 105.160 180.870 105.440 ;
        RECT 181.430 105.160 184.790 105.440 ;
        RECT 187.870 105.160 188.430 105.440 ;
        RECT 193.330 105.300 193.750 105.440 ;
        RECT 176.950 104.880 180.590 105.160 ;
        RECT 181.710 104.880 185.070 105.160 ;
        RECT 187.870 104.880 188.710 105.160 ;
        RECT 169.950 102.080 170.510 104.880 ;
        RECT 176.670 104.600 180.590 104.880 ;
        RECT 181.990 104.600 185.350 104.880 ;
        RECT 188.150 104.600 188.710 104.880 ;
        RECT 193.470 104.600 193.750 105.300 ;
        RECT 197.670 104.880 198.230 105.440 ;
        RECT 199.070 105.160 199.910 105.440 ;
        RECT 198.790 104.880 199.630 105.160 ;
        RECT 201.590 104.880 202.150 105.580 ;
        RECT 197.390 104.740 197.810 104.880 ;
        RECT 197.390 104.600 197.670 104.740 ;
        RECT 198.510 104.600 199.350 104.880 ;
        RECT 201.870 104.600 202.150 104.880 ;
        RECT 202.430 105.440 204.110 105.720 ;
        RECT 206.630 105.580 207.330 105.720 ;
        RECT 209.430 105.580 210.690 105.720 ;
        RECT 206.630 105.440 207.190 105.580 ;
        RECT 209.430 105.440 210.550 105.580 ;
        RECT 211.950 105.440 212.510 105.720 ;
        RECT 202.430 105.160 202.990 105.440 ;
        RECT 206.630 105.160 206.910 105.440 ;
        RECT 208.030 105.300 209.570 105.440 ;
        RECT 208.030 105.160 209.430 105.300 ;
        RECT 211.390 105.160 212.510 105.440 ;
        RECT 202.430 104.600 202.710 105.160 ;
        RECT 206.350 105.020 208.170 105.160 ;
        RECT 210.270 105.020 211.530 105.160 ;
        RECT 206.350 104.880 206.630 105.020 ;
        RECT 206.910 104.880 208.030 105.020 ;
        RECT 210.270 104.880 211.390 105.020 ;
        RECT 212.230 104.880 212.510 105.160 ;
        RECT 205.790 104.740 207.050 104.880 ;
        RECT 208.870 104.740 210.410 104.880 ;
        RECT 212.370 104.740 212.790 104.880 ;
        RECT 205.790 104.600 206.910 104.740 ;
        RECT 208.870 104.600 210.270 104.740 ;
        RECT 176.670 104.320 180.870 104.600 ;
        RECT 182.270 104.320 185.630 104.600 ;
        RECT 188.150 104.320 188.990 104.600 ;
        RECT 193.610 104.460 194.030 104.600 ;
        RECT 176.390 104.040 181.150 104.320 ;
        RECT 182.550 104.040 185.910 104.320 ;
        RECT 188.430 104.040 188.990 104.320 ;
        RECT 176.110 103.760 181.430 104.040 ;
        RECT 176.110 103.480 181.710 103.760 ;
        RECT 182.830 103.480 186.190 104.040 ;
        RECT 188.430 103.760 189.270 104.040 ;
        RECT 188.710 103.480 189.270 103.760 ;
        RECT 193.750 103.760 194.030 104.460 ;
        RECT 197.110 104.460 197.530 104.600 ;
        RECT 197.110 104.320 197.390 104.460 ;
        RECT 198.230 104.320 199.070 104.600 ;
        RECT 201.590 104.320 202.990 104.600 ;
        RECT 196.550 104.180 197.250 104.320 ;
        RECT 196.550 104.040 197.110 104.180 ;
        RECT 197.950 104.040 198.790 104.320 ;
        RECT 201.310 104.040 202.150 104.320 ;
        RECT 202.710 104.040 202.990 104.320 ;
        RECT 206.070 104.040 206.350 104.600 ;
        RECT 207.750 104.460 209.010 104.600 ;
        RECT 207.750 104.320 208.870 104.460 ;
        RECT 206.630 104.180 207.890 104.320 ;
        RECT 206.630 104.040 207.750 104.180 ;
        RECT 212.510 104.040 212.790 104.740 ;
        RECT 213.630 104.040 213.910 106.000 ;
        RECT 219.230 105.720 219.510 106.280 ;
        RECT 225.110 106.000 227.070 106.280 ;
        RECT 229.310 106.000 230.150 106.280 ;
        RECT 233.510 106.000 234.350 106.280 ;
        RECT 235.190 106.000 236.030 106.280 ;
        RECT 240.790 106.000 245.830 106.280 ;
        RECT 225.390 105.720 227.350 106.000 ;
        RECT 229.590 105.720 230.430 106.000 ;
        RECT 233.790 105.720 235.750 106.000 ;
        RECT 239.950 105.720 243.030 106.000 ;
        RECT 243.590 105.720 244.990 106.000 ;
        RECT 219.230 105.440 219.790 105.720 ;
        RECT 225.950 105.440 226.510 105.720 ;
        RECT 226.790 105.440 227.630 105.720 ;
        RECT 229.870 105.440 230.710 105.720 ;
        RECT 234.070 105.440 235.190 105.720 ;
        RECT 237.430 105.440 242.750 105.720 ;
        RECT 243.870 105.440 244.150 105.720 ;
        RECT 219.510 104.880 219.790 105.440 ;
        RECT 226.790 105.160 227.910 105.440 ;
        RECT 230.150 105.160 230.710 105.440 ;
        RECT 234.350 105.160 235.190 105.440 ;
        RECT 237.150 105.160 242.470 105.440 ;
        RECT 226.230 104.880 228.190 105.160 ;
        RECT 230.430 104.880 230.990 105.160 ;
        RECT 233.790 104.880 234.630 105.160 ;
        RECT 235.050 105.020 235.470 105.160 ;
        RECT 235.190 104.880 235.470 105.020 ;
        RECT 236.870 104.880 242.470 105.160 ;
        RECT 258.710 104.880 311.630 105.440 ;
        RECT 219.230 104.320 219.790 104.880 ;
        RECT 225.950 104.600 228.470 104.880 ;
        RECT 230.430 104.600 231.270 104.880 ;
        RECT 233.230 104.600 234.350 104.880 ;
        RECT 235.190 104.600 236.030 104.880 ;
        RECT 236.590 104.600 241.910 104.880 ;
        RECT 258.430 104.600 311.630 104.880 ;
        RECT 196.270 103.760 196.830 104.040 ;
        RECT 197.670 103.760 198.510 104.040 ;
        RECT 201.030 103.760 201.870 104.040 ;
        RECT 202.710 103.760 203.270 104.040 ;
        RECT 205.790 103.900 206.770 104.040 ;
        RECT 205.790 103.760 206.630 103.900 ;
        RECT 213.630 103.760 214.190 104.040 ;
        RECT 219.230 103.760 219.510 104.320 ;
        RECT 225.950 104.040 228.750 104.600 ;
        RECT 222.030 103.760 222.590 104.040 ;
        RECT 225.670 103.760 229.030 104.040 ;
        RECT 193.750 103.480 194.310 103.760 ;
        RECT 195.990 103.480 196.550 103.760 ;
        RECT 197.390 103.480 198.230 103.760 ;
        RECT 200.750 103.480 201.590 103.760 ;
        RECT 175.830 103.200 181.990 103.480 ;
        RECT 183.110 103.200 186.470 103.480 ;
        RECT 188.710 103.200 189.550 103.480 ;
        RECT 175.550 102.920 179.470 103.200 ;
        RECT 179.750 102.920 182.270 103.200 ;
        RECT 183.390 102.920 186.750 103.200 ;
        RECT 175.550 102.640 179.190 102.920 ;
        RECT 180.030 102.640 182.550 102.920 ;
        RECT 183.670 102.640 186.750 102.920 ;
        RECT 188.990 102.640 189.550 103.200 ;
        RECT 197.110 103.200 197.950 103.480 ;
        RECT 200.470 103.200 201.590 103.480 ;
        RECT 202.710 103.480 203.830 103.760 ;
        RECT 202.710 103.200 204.110 103.480 ;
        RECT 197.110 102.920 197.670 103.200 ;
        RECT 200.190 102.920 201.870 103.200 ;
        RECT 202.710 102.920 204.390 103.200 ;
        RECT 196.830 102.640 197.670 102.920 ;
        RECT 199.910 102.640 200.750 102.920 ;
        RECT 201.030 102.640 201.870 102.920 ;
        RECT 175.270 102.360 178.910 102.640 ;
        RECT 180.310 102.360 182.830 102.640 ;
        RECT 183.670 102.360 187.030 102.640 ;
        RECT 188.990 102.360 189.830 102.640 ;
        RECT 196.830 102.360 197.390 102.640 ;
        RECT 199.910 102.360 200.470 102.640 ;
        RECT 151.470 101.520 155.670 102.080 ;
        RECT 156.790 101.800 159.030 102.080 ;
        RECT 168.830 101.800 170.510 102.080 ;
        RECT 174.990 102.080 178.910 102.360 ;
        RECT 180.590 102.080 182.830 102.360 ;
        RECT 183.950 102.080 187.310 102.360 ;
        RECT 174.990 101.800 178.630 102.080 ;
        RECT 180.870 101.800 183.110 102.080 ;
        RECT 184.230 101.800 187.310 102.080 ;
        RECT 189.270 102.080 189.830 102.360 ;
        RECT 196.550 102.080 197.110 102.360 ;
        RECT 199.630 102.080 200.470 102.360 ;
        RECT 201.310 102.080 201.870 102.640 ;
        RECT 202.990 102.640 204.670 102.920 ;
        RECT 206.070 102.640 206.350 103.480 ;
        RECT 212.790 102.640 213.070 103.760 ;
        RECT 213.910 103.480 214.190 103.760 ;
        RECT 218.950 103.620 219.370 103.760 ;
        RECT 218.950 103.480 219.230 103.620 ;
        RECT 221.470 103.480 222.310 103.760 ;
        RECT 225.390 103.480 229.310 103.760 ;
        RECT 230.710 103.480 231.270 104.600 ;
        RECT 232.670 104.320 233.790 104.600 ;
        RECT 234.910 104.320 241.070 104.600 ;
        RECT 258.430 104.320 311.350 104.600 ;
        RECT 232.390 104.040 233.510 104.320 ;
        RECT 234.350 104.040 239.950 104.320 ;
        RECT 258.150 104.040 311.350 104.320 ;
        RECT 231.830 103.760 233.230 104.040 ;
        RECT 233.790 103.760 235.470 104.040 ;
        RECT 236.310 103.760 239.670 104.040 ;
        RECT 258.150 103.760 311.070 104.040 ;
        RECT 231.550 103.480 235.190 103.760 ;
        RECT 236.030 103.480 239.110 103.760 ;
        RECT 258.150 103.480 310.790 103.760 ;
        RECT 214.050 103.340 214.470 103.480 ;
        RECT 214.190 103.200 214.470 103.340 ;
        RECT 218.670 103.200 219.230 103.480 ;
        RECT 220.910 103.200 221.750 103.480 ;
        RECT 225.390 103.200 229.870 103.480 ;
        RECT 230.150 103.200 234.630 103.480 ;
        RECT 236.030 103.200 238.830 103.480 ;
        RECT 257.870 103.200 310.790 103.480 ;
        RECT 214.190 102.920 214.750 103.200 ;
        RECT 218.390 102.920 218.950 103.200 ;
        RECT 220.070 103.060 221.050 103.200 ;
        RECT 220.070 102.920 220.910 103.060 ;
        RECT 225.390 102.920 234.350 103.200 ;
        RECT 236.030 102.920 238.270 103.200 ;
        RECT 214.470 102.640 215.030 102.920 ;
        RECT 218.110 102.640 218.670 102.920 ;
        RECT 219.230 102.640 220.350 102.920 ;
        RECT 225.950 102.640 228.750 102.920 ;
        RECT 229.590 102.640 233.790 102.920 ;
        RECT 202.990 102.360 205.230 102.640 ;
        RECT 214.750 102.360 215.590 102.640 ;
        RECT 217.550 102.360 219.510 102.640 ;
        RECT 226.510 102.360 228.750 102.640 ;
        RECT 230.290 102.500 234.070 102.640 ;
        RECT 230.430 102.360 234.070 102.500 ;
        RECT 235.750 102.360 237.990 102.920 ;
        RECT 202.990 102.080 205.510 102.360 ;
        RECT 156.510 101.520 158.750 101.800 ;
        RECT 167.990 101.520 171.910 101.800 ;
        RECT 151.190 101.240 155.390 101.520 ;
        RECT 156.510 101.240 158.470 101.520 ;
        RECT 166.870 101.240 173.030 101.520 ;
        RECT 174.710 101.240 178.350 101.800 ;
        RECT 181.150 101.520 183.390 101.800 ;
        RECT 184.230 101.520 187.590 101.800 ;
        RECT 189.270 101.520 190.110 102.080 ;
        RECT 181.430 101.240 183.390 101.520 ;
        RECT 184.510 101.240 187.590 101.520 ;
        RECT 151.190 100.960 155.110 101.240 ;
        RECT 156.230 100.960 158.470 101.240 ;
        RECT 166.310 100.960 168.270 101.240 ;
        RECT 171.630 100.960 173.590 101.240 ;
        RECT 174.430 100.960 178.070 101.240 ;
        RECT 181.430 100.960 183.670 101.240 ;
        RECT 150.910 100.680 155.110 100.960 ;
        RECT 155.950 100.680 158.190 100.960 ;
        RECT 165.750 100.680 167.430 100.960 ;
        RECT 172.470 100.680 178.070 100.960 ;
        RECT 181.710 100.680 183.950 100.960 ;
        RECT 184.790 100.680 187.870 101.240 ;
        RECT 189.550 100.960 190.110 101.520 ;
        RECT 196.270 101.800 197.110 102.080 ;
        RECT 199.350 101.800 200.190 102.080 ;
        RECT 196.270 101.240 196.830 101.800 ;
        RECT 199.350 101.520 200.470 101.800 ;
        RECT 201.310 101.520 202.150 102.080 ;
        RECT 202.990 101.800 203.270 102.080 ;
        RECT 203.830 101.800 205.790 102.080 ;
        RECT 203.130 101.660 203.550 101.800 ;
        RECT 195.990 100.960 196.830 101.240 ;
        RECT 199.070 101.240 200.470 101.520 ;
        RECT 189.550 100.680 190.390 100.960 ;
        RECT 150.910 100.120 154.830 100.680 ;
        RECT 155.950 100.400 157.910 100.680 ;
        RECT 165.190 100.400 166.590 100.680 ;
        RECT 173.310 100.400 177.790 100.680 ;
        RECT 181.990 100.400 183.950 100.680 ;
        RECT 155.670 100.120 157.910 100.400 ;
        RECT 164.630 100.120 166.030 100.400 ;
        RECT 173.870 100.120 177.510 100.400 ;
        RECT 150.630 99.560 154.550 100.120 ;
        RECT 155.670 99.840 157.630 100.120 ;
        RECT 164.350 99.840 165.470 100.120 ;
        RECT 173.590 99.840 177.510 100.120 ;
        RECT 181.990 99.840 184.230 100.400 ;
        RECT 185.070 100.120 188.150 100.680 ;
        RECT 155.390 99.560 157.630 99.840 ;
        RECT 164.070 99.560 165.190 99.840 ;
        RECT 173.590 99.560 177.230 99.840 ;
        RECT 181.990 99.560 184.510 99.840 ;
        RECT 185.350 99.560 188.430 100.120 ;
        RECT 189.830 99.840 190.390 100.680 ;
        RECT 195.990 100.400 196.550 100.960 ;
        RECT 199.070 100.680 199.630 101.240 ;
        RECT 199.910 100.680 200.470 101.240 ;
        RECT 201.590 100.960 202.150 101.520 ;
        RECT 203.270 100.960 203.550 101.660 ;
        RECT 204.390 101.520 206.070 101.800 ;
        RECT 204.670 101.240 206.070 101.520 ;
        RECT 206.350 101.240 206.630 102.360 ;
        RECT 212.790 101.520 213.070 102.360 ;
        RECT 215.310 102.080 218.670 102.360 ;
        RECT 226.790 102.080 228.750 102.360 ;
        RECT 230.150 102.080 234.630 102.360 ;
        RECT 235.470 102.080 237.710 102.360 ;
        RECT 245.550 102.080 249.750 102.360 ;
        RECT 216.150 101.800 217.830 102.080 ;
        RECT 222.590 101.800 223.710 102.080 ;
        RECT 227.350 101.800 229.310 102.080 ;
        RECT 230.150 101.800 237.430 102.080 ;
        RECT 244.710 101.940 245.690 102.080 ;
        RECT 249.610 101.940 250.030 102.080 ;
        RECT 244.710 101.800 245.550 101.940 ;
        RECT 215.310 101.520 216.990 101.800 ;
        RECT 222.310 101.520 223.710 101.800 ;
        RECT 227.630 101.520 232.110 101.800 ;
        RECT 232.250 101.660 237.430 101.800 ;
        RECT 212.510 101.380 212.930 101.520 ;
        RECT 212.510 101.240 212.790 101.380 ;
        RECT 214.470 101.240 216.150 101.520 ;
        RECT 195.710 100.120 196.550 100.400 ;
        RECT 189.830 99.560 190.670 99.840 ;
        RECT 150.350 98.720 154.270 99.560 ;
        RECT 155.390 99.280 157.350 99.560 ;
        RECT 163.790 99.280 164.630 99.560 ;
        RECT 173.310 99.280 176.950 99.560 ;
        RECT 155.110 98.720 157.630 99.280 ;
        RECT 163.510 99.000 164.350 99.280 ;
        RECT 173.030 99.000 176.950 99.280 ;
        RECT 181.710 99.280 184.510 99.560 ;
        RECT 181.710 99.000 184.790 99.280 ;
        RECT 163.230 98.720 164.070 99.000 ;
        RECT 173.030 98.720 177.230 99.000 ;
        RECT 181.430 98.720 184.790 99.000 ;
        RECT 185.630 99.000 188.710 99.560 ;
        RECT 185.630 98.720 188.990 99.000 ;
        RECT 150.350 98.440 153.990 98.720 ;
        RECT 155.110 98.440 157.910 98.720 ;
        RECT 162.950 98.440 163.790 98.720 ;
        RECT 168.550 98.440 171.350 98.720 ;
        RECT 172.750 98.440 177.790 98.720 ;
        RECT 181.150 98.440 184.790 98.720 ;
        RECT 150.070 97.880 153.990 98.440 ;
        RECT 154.830 98.160 157.910 98.440 ;
        RECT 162.670 98.160 163.510 98.440 ;
        RECT 167.710 98.160 170.230 98.440 ;
        RECT 170.510 98.160 172.190 98.440 ;
        RECT 172.470 98.160 178.910 98.440 ;
        RECT 180.870 98.160 185.070 98.440 ;
        RECT 154.830 97.880 158.190 98.160 ;
        RECT 150.070 97.320 153.710 97.880 ;
        RECT 154.830 97.600 158.470 97.880 ;
        RECT 162.390 97.600 163.230 98.160 ;
        RECT 167.150 97.880 168.270 98.160 ;
        RECT 166.590 97.600 167.430 97.880 ;
        RECT 149.790 97.040 153.710 97.320 ;
        RECT 154.550 97.320 158.750 97.600 ;
        RECT 162.110 97.320 162.950 97.600 ;
        RECT 166.310 97.320 167.430 97.600 ;
        RECT 154.550 97.040 159.030 97.320 ;
        RECT 162.110 97.040 162.670 97.320 ;
        RECT 166.030 97.040 167.430 97.320 ;
        RECT 168.830 97.320 169.950 98.160 ;
        RECT 171.630 97.600 176.110 98.160 ;
        RECT 176.390 97.880 178.910 98.160 ;
        RECT 180.590 97.880 185.070 98.160 ;
        RECT 185.910 98.160 188.990 98.720 ;
        RECT 190.110 98.160 190.670 99.560 ;
        RECT 195.710 98.160 196.270 100.120 ;
        RECT 198.790 99.560 199.350 100.680 ;
        RECT 199.910 100.120 200.750 100.680 ;
        RECT 201.590 100.400 202.430 100.960 ;
        RECT 203.270 100.680 203.830 100.960 ;
        RECT 200.190 99.560 200.750 100.120 ;
        RECT 201.870 100.120 202.430 100.400 ;
        RECT 203.550 100.120 203.830 100.680 ;
        RECT 204.950 100.120 206.070 101.240 ;
        RECT 206.490 101.100 206.910 101.240 ;
        RECT 206.630 100.680 206.910 101.100 ;
        RECT 212.230 101.100 212.650 101.240 ;
        RECT 212.230 100.960 212.510 101.100 ;
        RECT 213.350 100.960 215.030 101.240 ;
        RECT 211.950 100.680 214.190 100.960 ;
        RECT 206.770 100.540 207.190 100.680 ;
        RECT 206.910 100.400 207.190 100.540 ;
        RECT 210.830 100.400 213.070 100.680 ;
        RECT 207.050 100.260 207.750 100.400 ;
        RECT 207.190 100.120 207.750 100.260 ;
        RECT 209.430 100.120 211.950 100.400 ;
        RECT 201.870 99.560 202.710 100.120 ;
        RECT 203.550 99.840 204.670 100.120 ;
        RECT 204.950 99.840 206.350 100.120 ;
        RECT 206.910 99.840 210.550 100.120 ;
        RECT 203.550 99.560 209.430 99.840 ;
        RECT 209.990 99.560 212.790 99.840 ;
        RECT 198.510 98.720 199.070 99.560 ;
        RECT 200.190 99.280 201.030 99.560 ;
        RECT 200.470 98.720 201.030 99.280 ;
        RECT 202.150 99.000 202.710 99.560 ;
        RECT 203.830 99.280 206.910 99.560 ;
        RECT 209.150 99.280 213.350 99.560 ;
        RECT 203.830 99.000 204.110 99.280 ;
        RECT 208.590 99.000 213.910 99.280 ;
        RECT 185.910 97.880 189.270 98.160 ;
        RECT 176.670 97.600 178.910 97.880 ;
        RECT 180.030 97.600 185.070 97.880 ;
        RECT 186.190 97.600 189.270 97.880 ;
        RECT 190.110 97.600 190.950 98.160 ;
        RECT 195.710 97.880 196.550 98.160 ;
        RECT 171.350 97.320 175.830 97.600 ;
        RECT 176.950 97.320 179.190 97.600 ;
        RECT 179.470 97.320 185.350 97.600 ;
        RECT 149.790 95.920 153.430 97.040 ;
        RECT 154.550 96.760 157.070 97.040 ;
        RECT 157.630 96.760 159.870 97.040 ;
        RECT 161.830 96.760 162.670 97.040 ;
        RECT 165.750 96.760 167.710 97.040 ;
        RECT 168.830 96.760 170.230 97.320 ;
        RECT 171.350 97.040 175.550 97.320 ;
        RECT 176.670 97.040 185.350 97.320 ;
        RECT 186.190 97.320 189.550 97.600 ;
        RECT 186.190 97.040 189.830 97.320 ;
        RECT 171.070 96.760 175.550 97.040 ;
        RECT 176.390 96.760 185.350 97.040 ;
        RECT 154.550 96.480 157.910 96.760 ;
        RECT 158.470 96.480 160.710 96.760 ;
        RECT 161.830 96.480 162.390 96.760 ;
        RECT 165.470 96.480 166.030 96.760 ;
        RECT 166.310 96.480 167.990 96.760 ;
        RECT 168.830 96.480 175.270 96.760 ;
        RECT 149.510 95.640 153.430 95.920 ;
        RECT 154.270 96.200 158.750 96.480 ;
        RECT 159.310 96.200 162.390 96.480 ;
        RECT 165.190 96.200 165.750 96.480 ;
        RECT 166.590 96.340 168.970 96.480 ;
        RECT 166.590 96.200 168.830 96.340 ;
        RECT 171.070 96.200 175.270 96.480 ;
        RECT 176.110 96.480 181.710 96.760 ;
        RECT 182.830 96.480 185.350 96.760 ;
        RECT 186.470 96.760 190.110 97.040 ;
        RECT 190.390 96.760 190.950 97.600 ;
        RECT 195.990 97.320 196.550 97.880 ;
        RECT 198.790 97.600 199.350 98.720 ;
        RECT 200.470 98.160 201.310 98.720 ;
        RECT 202.150 98.440 202.990 99.000 ;
        RECT 203.830 98.720 204.390 99.000 ;
        RECT 208.310 98.720 214.470 99.000 ;
        RECT 200.750 97.880 201.310 98.160 ;
        RECT 202.430 98.160 202.990 98.440 ;
        RECT 204.110 98.160 204.390 98.720 ;
        RECT 208.030 98.440 214.750 98.720 ;
        RECT 207.750 98.160 215.030 98.440 ;
        RECT 198.790 97.320 199.630 97.600 ;
        RECT 200.750 97.320 201.590 97.880 ;
        RECT 202.430 97.600 203.270 98.160 ;
        RECT 204.110 97.880 204.670 98.160 ;
        RECT 207.470 97.880 215.310 98.160 ;
        RECT 195.990 96.760 196.830 97.320 ;
        RECT 199.070 97.040 199.630 97.320 ;
        RECT 201.030 97.040 201.590 97.320 ;
        RECT 202.710 97.320 203.270 97.600 ;
        RECT 204.390 97.320 204.670 97.880 ;
        RECT 207.190 97.600 210.270 97.880 ;
        RECT 207.190 97.320 207.750 97.600 ;
        RECT 199.070 96.760 199.910 97.040 ;
        RECT 176.110 96.200 180.870 96.480 ;
        RECT 154.270 95.920 159.590 96.200 ;
        RECT 160.150 95.920 162.110 96.200 ;
        RECT 154.270 95.640 160.430 95.920 ;
        RECT 160.990 95.640 162.110 95.920 ;
        RECT 164.910 95.640 165.470 96.200 ;
        RECT 166.870 95.920 168.270 96.200 ;
        RECT 167.150 95.640 167.710 95.920 ;
        RECT 171.070 95.640 174.990 96.200 ;
        RECT 175.830 95.920 180.310 96.200 ;
        RECT 183.670 95.920 185.630 96.480 ;
        RECT 175.550 95.640 179.750 95.920 ;
        RECT 149.510 90.040 153.150 95.640 ;
        RECT 154.270 95.360 157.350 95.640 ;
        RECT 158.750 95.360 162.110 95.640 ;
        RECT 164.630 95.360 165.470 95.640 ;
        RECT 166.870 95.360 167.430 95.640 ;
        RECT 170.790 95.360 179.470 95.640 ;
        RECT 154.270 95.080 156.510 95.360 ;
        RECT 159.590 95.080 161.830 95.360 ;
        RECT 153.990 94.520 155.950 95.080 ;
        RECT 160.710 94.800 161.830 95.080 ;
        RECT 160.990 94.520 161.830 94.800 ;
        RECT 164.350 95.080 166.030 95.360 ;
        RECT 166.870 95.080 167.150 95.360 ;
        RECT 170.510 95.080 174.430 95.360 ;
        RECT 174.990 95.080 179.470 95.360 ;
        RECT 183.950 95.080 185.630 95.920 ;
        RECT 186.470 95.640 190.950 96.760 ;
        RECT 196.270 96.200 197.110 96.760 ;
        RECT 199.350 96.200 199.910 96.760 ;
        RECT 201.030 96.480 201.870 97.040 ;
        RECT 202.710 96.760 203.550 97.320 ;
        RECT 204.390 97.040 204.950 97.320 ;
        RECT 201.310 96.200 201.870 96.480 ;
        RECT 202.990 96.480 203.550 96.760 ;
        RECT 204.670 96.480 204.950 97.040 ;
        RECT 206.910 97.040 207.750 97.320 ;
        RECT 208.310 97.320 209.710 97.600 ;
        RECT 208.310 97.040 209.430 97.320 ;
        RECT 206.910 96.760 209.150 97.040 ;
        RECT 206.630 96.480 208.870 96.760 ;
        RECT 196.550 95.640 197.390 96.200 ;
        RECT 199.630 95.640 200.190 96.200 ;
        RECT 201.310 95.640 202.150 96.200 ;
        RECT 202.990 95.920 203.830 96.480 ;
        RECT 204.810 96.340 205.230 96.480 ;
        RECT 164.350 94.940 167.010 95.080 ;
        RECT 164.350 94.520 166.870 94.940 ;
        RECT 170.510 94.800 179.750 95.080 ;
        RECT 170.230 94.520 179.750 94.800 ;
        RECT 183.950 94.520 185.910 95.080 ;
        RECT 153.990 91.160 155.670 94.520 ;
        RECT 160.990 91.160 161.550 94.520 ;
        RECT 164.350 94.240 166.590 94.520 ;
        RECT 164.070 93.400 164.630 94.240 ;
        RECT 165.470 93.960 166.590 94.240 ;
        RECT 169.950 93.960 179.750 94.520 ;
        RECT 164.070 92.840 164.350 93.400 ;
        RECT 166.030 92.840 166.310 93.960 ;
        RECT 169.670 93.680 179.750 93.960 ;
        RECT 169.390 93.400 179.750 93.680 ;
        RECT 169.390 93.120 173.310 93.400 ;
        RECT 173.590 93.120 179.750 93.400 ;
        RECT 164.070 91.720 166.310 92.840 ;
        RECT 169.110 92.840 173.030 93.120 ;
        RECT 169.110 92.560 172.750 92.840 ;
        RECT 168.830 92.280 172.750 92.560 ;
        RECT 168.550 92.000 172.470 92.280 ;
        RECT 173.590 92.000 173.870 93.120 ;
        RECT 174.430 92.840 179.750 93.120 ;
        RECT 174.710 92.280 179.750 92.840 ;
        RECT 174.990 92.000 179.750 92.280 ;
        RECT 168.550 91.720 172.190 92.000 ;
        RECT 164.070 91.440 164.630 91.720 ;
        RECT 166.170 91.580 166.590 91.720 ;
        RECT 164.350 91.160 164.630 91.440 ;
        RECT 166.310 91.160 166.590 91.580 ;
        RECT 168.270 91.440 172.190 91.720 ;
        RECT 173.310 91.720 174.710 92.000 ;
        RECT 175.270 91.720 179.750 92.000 ;
        RECT 173.310 91.440 179.750 91.720 ;
        RECT 153.990 90.600 155.950 91.160 ;
        RECT 160.990 90.880 161.830 91.160 ;
        RECT 149.510 89.760 153.430 90.040 ;
        RECT 149.790 88.640 153.430 89.760 ;
        RECT 154.270 89.760 155.950 90.600 ;
        RECT 161.270 90.320 161.830 90.880 ;
        RECT 164.350 90.600 164.910 91.160 ;
        RECT 166.450 91.020 166.870 91.160 ;
        RECT 166.590 90.880 166.870 91.020 ;
        RECT 167.990 90.880 171.910 91.440 ;
        RECT 173.310 91.160 175.550 91.440 ;
        RECT 175.830 91.160 179.750 91.440 ;
        RECT 184.230 91.160 185.910 94.520 ;
        RECT 173.030 90.880 175.550 91.160 ;
        RECT 176.390 90.880 179.750 91.160 ;
        RECT 166.030 90.600 166.870 90.880 ;
        RECT 167.710 90.600 171.630 90.880 ;
        RECT 173.030 90.600 173.310 90.880 ;
        RECT 174.150 90.600 175.550 90.880 ;
        RECT 176.950 90.600 179.470 90.880 ;
        RECT 183.950 90.600 185.910 91.160 ;
        RECT 164.630 90.320 164.910 90.600 ;
        RECT 165.750 90.320 167.150 90.600 ;
        RECT 161.270 89.760 162.110 90.320 ;
        RECT 164.630 90.040 165.190 90.320 ;
        RECT 165.470 90.040 167.430 90.320 ;
        RECT 167.710 90.040 171.350 90.600 ;
        RECT 172.750 90.460 173.170 90.600 ;
        RECT 172.750 90.320 173.030 90.460 ;
        RECT 172.470 90.040 173.030 90.320 ;
        RECT 174.710 90.040 175.270 90.600 ;
        RECT 178.070 90.320 178.910 90.600 ;
        RECT 154.270 89.200 156.230 89.760 ;
        RECT 161.550 89.480 162.110 89.760 ;
        RECT 164.910 89.760 167.150 90.040 ;
        RECT 167.290 89.900 171.070 90.040 ;
        RECT 167.430 89.760 171.070 89.900 ;
        RECT 171.910 89.760 173.310 90.040 ;
        RECT 164.910 89.480 166.870 89.760 ;
        RECT 167.710 89.480 170.790 89.760 ;
        RECT 171.630 89.480 173.590 89.760 ;
        RECT 174.430 89.480 174.990 90.040 ;
        RECT 177.790 89.760 178.630 90.320 ;
        RECT 183.950 89.760 185.630 90.600 ;
        RECT 186.750 90.040 190.390 95.640 ;
        RECT 190.670 95.360 190.950 95.640 ;
        RECT 196.830 95.360 197.390 95.640 ;
        RECT 196.830 95.080 197.670 95.360 ;
        RECT 199.910 95.080 200.470 95.640 ;
        RECT 201.590 95.360 202.150 95.640 ;
        RECT 203.270 95.640 203.830 95.920 ;
        RECT 204.950 95.920 205.230 96.340 ;
        RECT 206.630 96.200 209.430 96.480 ;
        RECT 206.630 95.920 209.990 96.200 ;
        RECT 204.950 95.640 205.510 95.920 ;
        RECT 206.630 95.640 208.590 95.920 ;
        RECT 209.150 95.640 210.270 95.920 ;
        RECT 211.110 95.640 211.670 97.880 ;
        RECT 212.510 97.600 215.310 97.880 ;
        RECT 213.070 97.320 214.470 97.600 ;
        RECT 214.750 97.320 215.590 97.600 ;
        RECT 213.350 97.040 214.470 97.320 ;
        RECT 215.030 97.040 215.590 97.320 ;
        RECT 213.630 96.760 215.870 97.040 ;
        RECT 213.350 96.480 215.870 96.760 ;
        RECT 213.070 96.200 216.150 96.480 ;
        RECT 212.510 95.920 213.910 96.200 ;
        RECT 212.230 95.640 213.350 95.920 ;
        RECT 203.270 95.360 204.110 95.640 ;
        RECT 201.590 95.080 202.430 95.360 ;
        RECT 197.110 94.800 197.670 95.080 ;
        RECT 200.190 94.800 200.750 95.080 ;
        RECT 201.870 94.800 202.430 95.080 ;
        RECT 203.550 95.080 204.110 95.360 ;
        RECT 205.230 95.080 205.510 95.640 ;
        RECT 203.550 94.800 204.390 95.080 ;
        RECT 205.370 94.940 205.790 95.080 ;
        RECT 197.110 94.520 197.950 94.800 ;
        RECT 200.190 94.520 201.030 94.800 ;
        RECT 197.390 94.240 197.950 94.520 ;
        RECT 200.470 94.240 201.030 94.520 ;
        RECT 201.870 94.240 202.710 94.800 ;
        RECT 203.830 94.520 204.390 94.800 ;
        RECT 205.510 94.520 205.790 94.940 ;
        RECT 206.350 94.520 208.310 95.640 ;
        RECT 209.710 95.360 210.830 95.640 ;
        RECT 211.110 95.360 213.070 95.640 ;
        RECT 209.990 95.080 212.510 95.360 ;
        RECT 210.550 94.520 212.230 95.080 ;
        RECT 197.390 93.960 198.230 94.240 ;
        RECT 200.470 93.960 201.310 94.240 ;
        RECT 197.670 93.680 198.230 93.960 ;
        RECT 200.750 93.680 201.310 93.960 ;
        RECT 202.150 93.680 202.990 94.240 ;
        RECT 203.830 93.960 204.670 94.520 ;
        RECT 205.650 94.380 206.070 94.520 ;
        RECT 205.790 94.240 206.070 94.380 ;
        RECT 206.350 94.240 208.590 94.520 ;
        RECT 209.990 94.240 212.790 94.520 ;
        RECT 205.790 93.960 208.590 94.240 ;
        RECT 209.710 93.960 210.830 94.240 ;
        RECT 204.110 93.680 204.950 93.960 ;
        RECT 206.070 93.680 208.590 93.960 ;
        RECT 209.150 93.680 210.550 93.960 ;
        RECT 197.670 93.400 198.510 93.680 ;
        RECT 200.750 93.400 201.590 93.680 ;
        RECT 197.950 93.120 198.790 93.400 ;
        RECT 201.030 93.120 201.590 93.400 ;
        RECT 202.430 93.400 202.990 93.680 ;
        RECT 204.390 93.400 204.950 93.680 ;
        RECT 206.210 93.540 209.990 93.680 ;
        RECT 206.350 93.400 209.990 93.540 ;
        RECT 202.430 93.120 203.270 93.400 ;
        RECT 204.390 93.120 205.230 93.400 ;
        RECT 206.350 93.120 209.710 93.400 ;
        RECT 198.230 92.840 198.790 93.120 ;
        RECT 201.310 92.840 201.870 93.120 ;
        RECT 198.230 92.560 199.070 92.840 ;
        RECT 201.310 92.560 202.150 92.840 ;
        RECT 202.710 92.560 203.550 93.120 ;
        RECT 204.670 92.840 205.230 93.120 ;
        RECT 206.630 92.840 208.030 93.120 ;
        RECT 208.310 92.840 209.150 93.120 ;
        RECT 204.670 92.560 205.510 92.840 ;
        RECT 206.910 92.560 207.750 92.840 ;
        RECT 208.310 92.560 209.430 92.840 ;
        RECT 198.510 92.280 199.070 92.560 ;
        RECT 201.590 92.280 202.150 92.560 ;
        RECT 198.510 92.000 199.350 92.280 ;
        RECT 201.590 92.000 202.430 92.280 ;
        RECT 202.990 92.000 203.830 92.560 ;
        RECT 204.950 92.280 205.790 92.560 ;
        RECT 206.910 92.280 209.990 92.560 ;
        RECT 205.230 92.000 206.070 92.280 ;
        RECT 207.190 92.000 210.830 92.280 ;
        RECT 211.110 92.000 211.670 94.240 ;
        RECT 211.950 93.960 213.070 94.240 ;
        RECT 214.190 93.960 216.150 96.200 ;
        RECT 222.310 95.920 222.870 101.520 ;
        RECT 223.150 101.240 223.710 101.520 ;
        RECT 227.910 101.240 231.550 101.520 ;
        RECT 232.390 101.240 237.430 101.660 ;
        RECT 244.150 101.660 244.850 101.800 ;
        RECT 244.150 101.520 244.710 101.660 ;
        RECT 248.630 101.520 249.190 101.800 ;
        RECT 223.150 100.960 223.990 101.240 ;
        RECT 228.190 100.960 231.270 101.240 ;
        RECT 223.150 100.680 225.110 100.960 ;
        RECT 228.470 100.680 230.710 100.960 ;
        RECT 232.110 100.680 235.750 101.240 ;
        RECT 236.590 100.960 237.430 101.240 ;
        RECT 243.870 101.380 244.290 101.520 ;
        RECT 247.790 101.380 248.770 101.520 ;
        RECT 237.150 100.680 237.990 100.960 ;
        RECT 243.870 100.680 244.150 101.380 ;
        RECT 247.790 101.240 248.630 101.380 ;
        RECT 249.750 101.240 250.030 101.940 ;
        RECT 244.430 100.960 247.510 101.240 ;
        RECT 249.750 100.960 253.110 101.240 ;
        RECT 249.470 100.680 255.070 100.960 ;
        RECT 223.150 100.400 225.950 100.680 ;
        RECT 223.150 100.120 226.790 100.400 ;
        RECT 223.150 99.840 227.350 100.120 ;
        RECT 228.750 99.840 230.430 100.680 ;
        RECT 231.830 100.400 236.590 100.680 ;
        RECT 237.850 100.540 238.550 100.680 ;
        RECT 237.990 100.400 238.550 100.540 ;
        RECT 243.310 100.400 244.150 100.680 ;
        RECT 248.910 100.400 250.030 100.680 ;
        RECT 252.270 100.400 256.470 100.680 ;
        RECT 231.830 100.120 237.430 100.400 ;
        RECT 238.410 100.260 238.830 100.400 ;
        RECT 238.550 100.120 238.830 100.260 ;
        RECT 242.470 100.120 244.150 100.400 ;
        RECT 248.350 100.120 250.030 100.400 ;
        RECT 254.510 100.120 257.590 100.400 ;
        RECT 223.150 99.560 227.630 99.840 ;
        RECT 223.150 99.280 227.910 99.560 ;
        RECT 228.470 99.280 230.710 99.840 ;
        RECT 231.550 99.560 238.270 100.120 ;
        RECT 241.910 99.840 245.270 100.120 ;
        RECT 246.950 99.840 250.310 100.120 ;
        RECT 255.910 99.840 258.710 100.120 ;
        RECT 241.350 99.560 243.030 99.840 ;
        RECT 243.310 99.560 253.110 99.840 ;
        RECT 257.030 99.560 259.550 99.840 ;
        RECT 231.270 99.280 238.270 99.560 ;
        RECT 240.790 99.280 242.190 99.560 ;
        RECT 243.310 99.280 255.070 99.560 ;
        RECT 258.150 99.280 260.390 99.560 ;
        RECT 223.150 99.000 230.150 99.280 ;
        RECT 231.270 99.000 237.990 99.280 ;
        RECT 240.230 99.000 241.630 99.280 ;
        RECT 243.310 99.000 256.470 99.280 ;
        RECT 258.990 99.000 260.950 99.280 ;
        RECT 223.150 98.720 228.750 99.000 ;
        RECT 230.710 98.720 237.990 99.000 ;
        RECT 239.950 98.720 241.070 99.000 ;
        RECT 243.310 98.720 250.590 99.000 ;
        RECT 253.950 98.720 257.590 99.000 ;
        RECT 259.830 98.720 261.790 99.000 ;
        RECT 223.150 98.440 227.350 98.720 ;
        RECT 229.310 98.440 237.710 98.720 ;
        RECT 239.390 98.440 240.510 98.720 ;
        RECT 242.750 98.440 250.870 98.720 ;
        RECT 255.630 98.440 258.710 98.720 ;
        RECT 260.390 98.440 262.350 98.720 ;
        RECT 223.150 98.160 225.950 98.440 ;
        RECT 227.910 98.160 237.710 98.440 ;
        RECT 239.110 98.160 240.230 98.440 ;
        RECT 242.190 98.160 250.870 98.440 ;
        RECT 256.750 98.160 259.550 98.440 ;
        RECT 261.230 98.160 262.910 98.440 ;
        RECT 223.150 97.880 224.830 98.160 ;
        RECT 226.510 97.880 237.430 98.160 ;
        RECT 238.830 97.880 239.950 98.160 ;
        RECT 241.350 97.880 243.030 98.160 ;
        RECT 243.590 97.880 250.870 98.160 ;
        RECT 257.870 97.880 260.110 98.160 ;
        RECT 261.790 97.880 263.470 98.160 ;
        RECT 223.150 97.600 224.270 97.880 ;
        RECT 225.110 97.600 236.870 97.880 ;
        RECT 238.550 97.600 239.670 97.880 ;
        RECT 240.790 97.600 242.190 97.880 ;
        RECT 223.150 95.920 223.990 97.600 ;
        RECT 224.550 97.320 229.030 97.600 ;
        RECT 224.270 96.200 224.830 97.320 ;
        RECT 225.670 97.040 227.630 97.320 ;
        RECT 225.670 96.760 226.510 97.040 ;
        RECT 228.190 96.760 229.870 97.040 ;
        RECT 230.150 96.760 235.470 97.600 ;
        RECT 238.270 97.320 239.390 97.600 ;
        RECT 240.510 97.320 241.350 97.600 ;
        RECT 238.270 97.040 239.110 97.320 ;
        RECT 239.950 97.040 240.790 97.320 ;
        RECT 243.870 97.040 251.150 97.880 ;
        RECT 258.990 97.600 260.950 97.880 ;
        RECT 262.350 97.600 263.750 97.880 ;
        RECT 259.830 97.320 261.510 97.600 ;
        RECT 262.910 97.320 264.310 97.600 ;
        RECT 260.670 97.040 262.350 97.320 ;
        RECT 263.470 97.040 264.590 97.320 ;
        RECT 237.990 96.760 238.830 97.040 ;
        RECT 239.670 96.760 240.230 97.040 ;
        RECT 244.150 96.760 251.150 97.040 ;
        RECT 261.230 96.760 262.350 97.040 ;
        RECT 263.750 96.760 265.150 97.040 ;
        RECT 225.670 96.480 226.230 96.760 ;
        RECT 226.790 96.480 235.470 96.760 ;
        RECT 236.030 96.480 238.550 96.760 ;
        RECT 225.670 96.200 225.950 96.480 ;
        RECT 226.510 96.200 238.550 96.480 ;
        RECT 244.150 96.200 251.430 96.760 ;
        RECT 264.310 96.480 265.430 96.760 ;
        RECT 264.590 96.200 265.990 96.480 ;
        RECT 224.550 95.920 225.950 96.200 ;
        RECT 222.310 95.360 222.590 95.920 ;
        RECT 212.510 93.680 213.630 93.960 ;
        RECT 213.910 93.680 216.150 93.960 ;
        RECT 212.790 93.400 215.870 93.680 ;
        RECT 213.350 92.840 215.870 93.400 ;
        RECT 213.070 92.560 215.590 92.840 ;
        RECT 212.790 92.280 214.190 92.560 ;
        RECT 214.750 92.280 215.590 92.560 ;
        RECT 222.030 92.280 222.590 95.360 ;
        RECT 223.150 95.360 224.270 95.920 ;
        RECT 224.830 95.360 225.950 95.920 ;
        RECT 226.230 95.640 238.270 96.200 ;
        RECT 226.510 95.360 238.270 95.640 ;
        RECT 244.430 95.920 251.430 96.200 ;
        RECT 265.150 95.920 266.270 96.200 ;
        RECT 244.430 95.640 251.710 95.920 ;
        RECT 265.430 95.640 266.550 95.920 ;
        RECT 244.430 95.360 246.390 95.640 ;
        RECT 250.310 95.360 251.710 95.640 ;
        RECT 265.710 95.360 266.830 95.640 ;
        RECT 223.150 95.080 224.550 95.360 ;
        RECT 225.110 95.080 226.230 95.360 ;
        RECT 223.150 94.800 224.830 95.080 ;
        RECT 225.390 94.800 226.230 95.080 ;
        RECT 226.790 94.800 237.990 95.360 ;
        RECT 244.430 95.080 246.110 95.360 ;
        RECT 250.590 95.080 251.710 95.360 ;
        RECT 265.990 95.080 267.110 95.360 ;
        RECT 223.150 94.520 225.110 94.800 ;
        RECT 225.670 94.520 226.510 94.800 ;
        RECT 227.070 94.520 237.990 94.800 ;
        RECT 223.150 93.680 223.990 94.520 ;
        RECT 224.270 94.240 225.390 94.520 ;
        RECT 225.950 94.240 226.790 94.520 ;
        RECT 227.350 94.240 234.910 94.520 ;
        RECT 224.270 93.960 225.670 94.240 ;
        RECT 222.870 93.400 223.990 93.680 ;
        RECT 224.550 93.680 225.670 93.960 ;
        RECT 226.230 93.960 227.070 94.240 ;
        RECT 226.230 93.680 227.350 93.960 ;
        RECT 227.630 93.680 234.630 94.240 ;
        RECT 224.550 93.400 225.950 93.680 ;
        RECT 226.510 93.400 227.350 93.680 ;
        RECT 227.910 93.400 234.350 93.680 ;
        RECT 236.590 93.400 237.990 94.520 ;
        RECT 244.710 94.800 246.110 95.080 ;
        RECT 246.670 94.800 250.030 95.080 ;
        RECT 250.590 94.800 251.990 95.080 ;
        RECT 266.270 94.800 267.390 95.080 ;
        RECT 244.710 94.240 246.390 94.800 ;
        RECT 246.670 94.520 249.750 94.800 ;
        RECT 246.950 94.240 249.750 94.520 ;
        RECT 250.310 94.240 251.990 94.800 ;
        RECT 266.550 94.520 267.670 94.800 ;
        RECT 266.830 94.240 267.950 94.520 ;
        RECT 244.990 93.680 246.670 94.240 ;
        RECT 246.950 93.960 249.470 94.240 ;
        RECT 250.030 93.960 252.270 94.240 ;
        RECT 267.110 93.960 268.230 94.240 ;
        RECT 247.230 93.680 249.470 93.960 ;
        RECT 244.990 93.400 246.950 93.680 ;
        RECT 222.870 92.280 224.270 93.400 ;
        RECT 211.950 92.000 215.310 92.280 ;
        RECT 222.310 92.000 224.270 92.280 ;
        RECT 198.790 91.720 199.350 92.000 ;
        RECT 201.870 91.720 202.430 92.000 ;
        RECT 203.270 91.720 204.110 92.000 ;
        RECT 205.230 91.720 206.350 92.000 ;
        RECT 207.470 91.720 215.030 92.000 ;
        RECT 222.590 91.720 224.270 92.000 ;
        RECT 198.790 91.440 199.630 91.720 ;
        RECT 199.070 91.160 199.630 91.440 ;
        RECT 202.150 91.440 202.710 91.720 ;
        RECT 203.550 91.440 204.390 91.720 ;
        RECT 205.510 91.440 206.630 91.720 ;
        RECT 207.750 91.440 214.750 91.720 ;
        RECT 202.150 91.160 202.990 91.440 ;
        RECT 199.070 90.880 199.910 91.160 ;
        RECT 202.430 90.880 202.990 91.160 ;
        RECT 203.830 91.160 204.390 91.440 ;
        RECT 205.790 91.160 206.910 91.440 ;
        RECT 208.030 91.160 214.470 91.440 ;
        RECT 223.150 91.160 224.270 91.720 ;
        RECT 224.550 93.120 226.230 93.400 ;
        RECT 226.790 93.120 227.630 93.400 ;
        RECT 228.190 93.120 234.350 93.400 ;
        RECT 224.550 92.840 226.510 93.120 ;
        RECT 227.070 92.840 234.070 93.120 ;
        RECT 224.550 92.560 226.790 92.840 ;
        RECT 227.350 92.560 233.790 92.840 ;
        RECT 224.550 92.000 227.070 92.560 ;
        RECT 227.630 92.280 233.790 92.560 ;
        RECT 236.870 92.280 237.990 93.400 ;
        RECT 245.270 92.840 247.230 93.400 ;
        RECT 247.510 93.120 249.190 93.680 ;
        RECT 249.750 93.400 252.270 93.960 ;
        RECT 267.390 93.680 268.510 93.960 ;
        RECT 267.670 93.400 268.790 93.680 ;
        RECT 247.790 92.840 248.910 93.120 ;
        RECT 249.470 92.840 252.550 93.400 ;
        RECT 267.950 93.120 268.790 93.400 ;
        RECT 268.230 92.840 269.070 93.120 ;
        RECT 245.270 92.280 247.510 92.840 ;
        RECT 247.790 92.560 248.630 92.840 ;
        RECT 249.190 92.560 252.550 92.840 ;
        RECT 248.070 92.280 248.630 92.560 ;
        RECT 248.910 92.280 252.550 92.560 ;
        RECT 268.510 92.560 269.350 92.840 ;
        RECT 268.510 92.280 269.630 92.560 ;
        RECT 227.630 92.000 233.510 92.280 ;
        RECT 224.550 91.440 233.510 92.000 ;
        RECT 237.150 92.000 237.990 92.280 ;
        RECT 237.150 91.440 238.270 92.000 ;
        RECT 245.550 91.720 247.790 92.280 ;
        RECT 248.910 92.000 252.830 92.280 ;
        RECT 268.790 92.000 269.630 92.280 ;
        RECT 248.630 91.720 252.830 92.000 ;
        RECT 245.550 91.440 252.830 91.720 ;
        RECT 269.070 91.440 269.910 92.000 ;
        RECT 224.550 91.160 226.510 91.440 ;
        RECT 226.930 91.300 233.790 91.440 ;
        RECT 227.070 91.160 233.790 91.300 ;
        RECT 203.830 90.880 204.670 91.160 ;
        RECT 206.070 90.880 207.190 91.160 ;
        RECT 208.590 90.880 214.190 91.160 ;
        RECT 223.430 90.880 225.950 91.160 ;
        RECT 227.070 90.880 234.350 91.160 ;
        RECT 237.430 90.880 238.270 91.440 ;
        RECT 199.350 90.600 200.190 90.880 ;
        RECT 202.430 90.600 203.270 90.880 ;
        RECT 204.110 90.600 204.950 90.880 ;
        RECT 206.630 90.600 207.470 90.880 ;
        RECT 208.870 90.600 213.630 90.880 ;
        RECT 223.430 90.600 225.390 90.880 ;
        RECT 226.790 90.600 234.910 90.880 ;
        RECT 199.630 90.320 200.190 90.600 ;
        RECT 202.710 90.320 203.270 90.600 ;
        RECT 204.390 90.320 205.230 90.600 ;
        RECT 206.910 90.320 208.030 90.600 ;
        RECT 209.710 90.320 213.070 90.600 ;
        RECT 226.790 90.320 235.190 90.600 ;
        RECT 237.430 90.320 238.550 90.880 ;
        RECT 245.830 90.600 253.110 91.440 ;
        RECT 269.350 90.880 270.190 91.440 ;
        RECT 199.630 90.040 200.470 90.320 ;
        RECT 177.790 89.480 178.350 89.760 ;
        RECT 161.550 89.200 162.390 89.480 ;
        RECT 165.190 89.200 166.310 89.480 ;
        RECT 167.990 89.200 170.790 89.480 ;
        RECT 171.070 89.340 171.770 89.480 ;
        RECT 171.070 89.200 171.630 89.340 ;
        RECT 172.190 89.200 173.590 89.480 ;
        RECT 174.150 89.200 174.710 89.480 ;
        RECT 177.510 89.200 178.350 89.480 ;
        RECT 183.670 89.200 185.630 89.760 ;
        RECT 186.470 89.760 190.390 90.040 ;
        RECT 199.910 89.760 200.470 90.040 ;
        RECT 202.990 90.040 203.550 90.320 ;
        RECT 204.670 90.040 205.510 90.320 ;
        RECT 207.470 90.040 208.590 90.320 ;
        RECT 210.830 90.040 211.950 90.320 ;
        RECT 226.510 90.040 235.750 90.320 ;
        RECT 237.710 90.040 238.550 90.320 ;
        RECT 202.990 89.760 203.830 90.040 ;
        RECT 204.950 89.760 206.070 90.040 ;
        RECT 207.750 89.760 209.150 90.040 ;
        RECT 226.510 89.760 236.310 90.040 ;
        RECT 154.550 88.640 156.230 89.200 ;
        RECT 161.830 88.920 162.390 89.200 ;
        RECT 165.470 88.920 166.030 89.200 ;
        RECT 167.710 89.060 171.210 89.200 ;
        RECT 161.830 88.640 162.670 88.920 ;
        RECT 165.750 88.640 166.310 88.920 ;
        RECT 167.710 88.640 171.070 89.060 ;
        RECT 172.190 88.920 174.430 89.200 ;
        RECT 177.510 88.920 178.070 89.200 ;
        RECT 172.470 88.640 174.150 88.920 ;
        RECT 177.230 88.640 178.070 88.920 ;
        RECT 183.670 88.640 185.350 89.200 ;
        RECT 186.470 88.640 190.110 89.760 ;
        RECT 199.910 89.480 200.750 89.760 ;
        RECT 203.270 89.480 203.830 89.760 ;
        RECT 205.230 89.480 206.350 89.760 ;
        RECT 208.310 89.480 209.990 89.760 ;
        RECT 226.230 89.480 236.870 89.760 ;
        RECT 237.710 89.480 238.830 90.040 ;
        RECT 246.110 89.760 253.390 90.600 ;
        RECT 269.630 90.320 270.470 90.880 ;
        RECT 269.910 89.760 270.750 90.320 ;
        RECT 246.110 89.480 253.670 89.760 ;
        RECT 200.190 89.200 200.750 89.480 ;
        RECT 203.550 89.200 204.110 89.480 ;
        RECT 205.510 89.200 206.910 89.480 ;
        RECT 209.150 89.200 211.110 89.480 ;
        RECT 226.230 89.200 232.390 89.480 ;
        RECT 232.950 89.200 237.150 89.480 ;
        RECT 237.710 89.200 239.110 89.480 ;
        RECT 200.470 88.920 201.030 89.200 ;
        RECT 203.550 88.920 204.390 89.200 ;
        RECT 206.070 88.920 207.190 89.200 ;
        RECT 209.990 88.920 211.950 89.200 ;
        RECT 200.470 88.640 201.310 88.920 ;
        RECT 203.830 88.640 204.390 88.920 ;
        RECT 206.350 88.640 208.030 88.920 ;
        RECT 211.390 88.640 211.950 88.920 ;
        RECT 225.950 88.640 232.110 89.200 ;
        RECT 233.510 88.920 239.110 89.200 ;
        RECT 233.790 88.640 239.390 88.920 ;
        RECT 246.390 88.640 253.670 89.480 ;
        RECT 149.790 88.360 153.710 88.640 ;
        RECT 150.070 87.800 153.710 88.360 ;
        RECT 154.550 88.080 156.510 88.640 ;
        RECT 162.110 88.360 162.670 88.640 ;
        RECT 166.030 88.360 166.590 88.640 ;
        RECT 162.110 88.080 162.950 88.360 ;
        RECT 166.310 88.080 167.150 88.360 ;
        RECT 167.430 88.080 168.830 88.640 ;
        RECT 154.830 87.800 156.510 88.080 ;
        RECT 162.390 87.800 163.230 88.080 ;
        RECT 166.590 87.800 168.550 88.080 ;
        RECT 169.950 87.800 171.350 88.640 ;
        RECT 172.750 88.360 173.870 88.640 ;
        RECT 177.230 88.360 177.790 88.640 ;
        RECT 172.750 88.080 173.590 88.360 ;
        RECT 176.950 88.080 177.790 88.360 ;
        RECT 183.390 88.080 185.350 88.640 ;
        RECT 186.190 88.360 190.110 88.640 ;
        RECT 200.750 88.360 201.310 88.640 ;
        RECT 172.470 87.800 173.310 88.080 ;
        RECT 176.670 87.800 177.510 88.080 ;
        RECT 183.390 87.800 185.070 88.080 ;
        RECT 186.190 87.800 189.830 88.360 ;
        RECT 200.750 88.080 201.590 88.360 ;
        RECT 204.110 88.080 204.670 88.640 ;
        RECT 206.910 88.360 208.590 88.640 ;
        RECT 207.470 88.080 209.430 88.360 ;
        RECT 225.670 88.080 231.830 88.640 ;
        RECT 234.350 88.360 239.670 88.640 ;
        RECT 234.910 88.080 239.950 88.360 ;
        RECT 201.030 87.800 201.590 88.080 ;
        RECT 204.390 87.800 204.950 88.080 ;
        RECT 208.310 87.800 210.550 88.080 ;
        RECT 225.390 87.800 231.830 88.080 ;
        RECT 235.470 87.800 240.510 88.080 ;
        RECT 246.670 87.800 253.950 88.640 ;
        RECT 150.070 87.240 153.990 87.800 ;
        RECT 154.830 87.240 156.790 87.800 ;
        RECT 162.670 87.520 163.230 87.800 ;
        RECT 167.150 87.520 168.550 87.800 ;
        RECT 170.230 87.520 171.350 87.800 ;
        RECT 171.630 87.520 172.750 87.800 ;
        RECT 176.670 87.520 177.230 87.800 ;
        RECT 162.670 87.240 163.510 87.520 ;
        RECT 167.710 87.240 169.670 87.520 ;
        RECT 169.950 87.240 172.190 87.520 ;
        RECT 176.390 87.240 177.230 87.520 ;
        RECT 183.110 87.240 185.070 87.800 ;
        RECT 185.910 87.240 189.830 87.800 ;
        RECT 201.310 87.520 201.870 87.800 ;
        RECT 201.310 87.240 202.150 87.520 ;
        RECT 204.670 87.240 205.230 87.800 ;
        RECT 209.150 87.520 211.390 87.800 ;
        RECT 210.270 87.240 211.390 87.520 ;
        RECT 225.110 87.240 231.550 87.800 ;
        RECT 236.030 87.520 240.790 87.800 ;
        RECT 236.310 87.240 241.350 87.520 ;
        RECT 150.350 86.960 153.990 87.240 ;
        RECT 150.350 86.120 154.270 86.960 ;
        RECT 155.110 86.680 157.070 87.240 ;
        RECT 162.950 86.960 163.790 87.240 ;
        RECT 168.830 86.960 171.070 87.240 ;
        RECT 176.110 86.960 176.950 87.240 ;
        RECT 163.230 86.680 164.070 86.960 ;
        RECT 175.830 86.680 176.670 86.960 ;
        RECT 182.830 86.680 184.790 87.240 ;
        RECT 185.910 86.960 189.550 87.240 ;
        RECT 201.590 86.960 202.150 87.240 ;
        RECT 204.950 86.960 205.510 87.240 ;
        RECT 155.110 86.400 157.350 86.680 ;
        RECT 163.510 86.400 164.350 86.680 ;
        RECT 175.550 86.400 176.390 86.680 ;
        RECT 155.390 86.120 157.350 86.400 ;
        RECT 163.790 86.120 164.630 86.400 ;
        RECT 175.270 86.120 176.670 86.400 ;
        RECT 182.550 86.120 184.510 86.680 ;
        RECT 185.630 86.400 189.550 86.960 ;
        RECT 201.870 86.680 202.430 86.960 ;
        RECT 201.870 86.400 202.710 86.680 ;
        RECT 205.230 86.400 205.790 86.960 ;
        RECT 224.830 86.680 231.270 87.240 ;
        RECT 236.310 86.960 241.910 87.240 ;
        RECT 246.950 86.960 254.230 87.800 ;
        RECT 224.550 86.400 231.270 86.680 ;
        RECT 236.030 86.680 242.750 86.960 ;
        RECT 246.950 86.680 254.510 86.960 ;
        RECT 236.030 86.400 243.590 86.680 ;
        RECT 150.630 85.560 154.550 86.120 ;
        RECT 155.390 85.840 157.630 86.120 ;
        RECT 155.670 85.560 157.630 85.840 ;
        RECT 164.070 85.840 165.190 86.120 ;
        RECT 174.710 85.840 176.950 86.120 ;
        RECT 182.270 85.840 184.510 86.120 ;
        RECT 185.350 86.120 189.550 86.400 ;
        RECT 202.150 86.120 202.710 86.400 ;
        RECT 205.510 86.120 206.070 86.400 ;
        RECT 224.550 86.120 230.990 86.400 ;
        RECT 164.070 85.560 165.470 85.840 ;
        RECT 174.430 85.560 177.230 85.840 ;
        RECT 182.270 85.560 184.230 85.840 ;
        RECT 185.350 85.560 189.270 86.120 ;
        RECT 202.430 85.840 202.990 86.120 ;
        RECT 202.430 85.560 203.270 85.840 ;
        RECT 224.270 85.560 230.990 86.120 ;
        RECT 236.030 85.840 237.150 86.400 ;
        RECT 150.910 85.000 154.830 85.560 ;
        RECT 155.670 85.280 157.910 85.560 ;
        RECT 164.070 85.280 166.030 85.560 ;
        RECT 173.870 85.280 174.990 85.560 ;
        RECT 175.270 85.280 177.230 85.560 ;
        RECT 181.990 85.280 184.230 85.560 ;
        RECT 155.950 85.000 157.910 85.280 ;
        RECT 163.790 85.000 166.590 85.280 ;
        RECT 173.310 85.000 174.710 85.280 ;
        RECT 175.550 85.000 177.510 85.280 ;
        RECT 181.990 85.000 183.950 85.280 ;
        RECT 185.070 85.000 188.990 85.560 ;
        RECT 202.710 85.280 203.270 85.560 ;
        RECT 150.910 84.720 155.110 85.000 ;
        RECT 155.950 84.720 158.190 85.000 ;
        RECT 151.190 84.440 155.110 84.720 ;
        RECT 156.230 84.440 158.470 84.720 ;
        RECT 163.510 84.440 165.470 85.000 ;
        RECT 165.750 84.720 167.430 85.000 ;
        RECT 172.470 84.720 174.150 85.000 ;
        RECT 175.550 84.720 177.790 85.000 ;
        RECT 181.710 84.720 183.950 85.000 ;
        RECT 184.790 84.720 188.990 85.000 ;
        RECT 202.990 84.720 203.550 85.280 ;
        RECT 223.990 85.000 230.710 85.560 ;
        RECT 223.710 84.720 230.710 85.000 ;
        RECT 235.750 85.000 237.150 85.840 ;
        RECT 237.710 86.120 245.270 86.400 ;
        RECT 247.230 86.120 254.510 86.680 ;
        RECT 267.390 86.120 269.350 86.400 ;
        RECT 237.710 85.840 254.790 86.120 ;
        RECT 261.790 85.840 269.350 86.120 ;
        RECT 237.710 85.560 269.070 85.840 ;
        RECT 237.710 85.280 264.310 85.560 ;
        RECT 237.990 85.000 239.950 85.280 ;
        RECT 240.510 85.000 256.750 85.280 ;
        RECT 166.310 84.440 168.550 84.720 ;
        RECT 171.350 84.440 173.590 84.720 ;
        RECT 175.830 84.440 178.070 84.720 ;
        RECT 181.430 84.440 183.670 84.720 ;
        RECT 184.790 84.440 188.710 84.720 ;
        RECT 203.270 84.440 203.830 84.720 ;
        RECT 223.710 84.440 230.430 84.720 ;
        RECT 151.190 84.160 155.390 84.440 ;
        RECT 151.470 83.600 155.670 84.160 ;
        RECT 156.510 83.880 158.750 84.440 ;
        RECT 163.230 84.160 165.190 84.440 ;
        RECT 167.150 84.160 172.750 84.440 ;
        RECT 176.110 84.160 178.350 84.440 ;
        RECT 162.950 83.880 164.910 84.160 ;
        RECT 167.990 83.880 171.910 84.160 ;
        RECT 176.390 83.880 178.630 84.160 ;
        RECT 181.150 83.880 183.390 84.440 ;
        RECT 184.510 84.160 188.710 84.440 ;
        RECT 156.790 83.600 159.030 83.880 ;
        RECT 162.670 83.600 164.910 83.880 ;
        RECT 176.390 83.600 178.910 83.880 ;
        RECT 180.870 83.600 183.110 83.880 ;
        RECT 184.230 83.600 188.430 84.160 ;
        RECT 203.550 83.880 204.110 84.440 ;
        RECT 223.430 83.880 230.430 84.440 ;
        RECT 235.750 83.880 237.430 85.000 ;
        RECT 237.990 84.160 240.230 85.000 ;
        RECT 241.070 84.720 257.310 85.000 ;
        RECT 241.630 84.440 258.710 84.720 ;
        RECT 242.190 84.160 258.990 84.440 ;
        RECT 238.270 83.880 240.230 84.160 ;
        RECT 242.470 83.880 259.550 84.160 ;
        RECT 151.750 83.320 155.950 83.600 ;
        RECT 157.070 83.320 159.310 83.600 ;
        RECT 162.670 83.320 164.630 83.600 ;
        RECT 176.670 83.320 180.030 83.600 ;
        RECT 180.590 83.320 182.830 83.600 ;
        RECT 183.950 83.320 188.150 83.600 ;
        RECT 223.150 83.320 230.150 83.880 ;
        RECT 151.750 83.040 156.230 83.320 ;
        RECT 157.070 83.040 159.590 83.320 ;
        RECT 162.110 83.040 164.350 83.320 ;
        RECT 152.030 82.760 156.230 83.040 ;
        RECT 157.350 82.760 159.870 83.040 ;
        RECT 161.550 82.760 164.350 83.040 ;
        RECT 176.950 83.040 182.830 83.320 ;
        RECT 183.670 83.040 188.150 83.320 ;
        RECT 222.870 83.040 230.150 83.320 ;
        RECT 236.030 83.040 237.710 83.880 ;
        RECT 238.270 83.040 240.510 83.880 ;
        RECT 243.030 83.600 259.830 83.880 ;
        RECT 243.590 83.320 260.110 83.600 ;
        RECT 243.590 83.040 260.390 83.320 ;
        RECT 176.950 82.760 182.550 83.040 ;
        RECT 183.670 82.760 187.870 83.040 ;
        RECT 222.870 82.760 229.310 83.040 ;
        RECT 236.030 82.760 237.990 83.040 ;
        RECT 152.030 82.480 156.510 82.760 ;
        RECT 157.630 82.480 164.070 82.760 ;
        RECT 176.950 82.480 182.270 82.760 ;
        RECT 183.390 82.480 187.870 82.760 ;
        RECT 222.590 82.480 228.190 82.760 ;
        RECT 152.310 82.200 156.790 82.480 ;
        RECT 157.910 82.200 164.070 82.480 ;
        RECT 177.230 82.200 181.990 82.480 ;
        RECT 183.110 82.200 187.590 82.480 ;
        RECT 222.590 82.200 227.350 82.480 ;
        RECT 152.590 81.920 157.070 82.200 ;
        RECT 158.190 81.920 163.790 82.200 ;
        RECT 177.230 81.920 181.710 82.200 ;
        RECT 182.830 81.920 187.310 82.200 ;
        RECT 152.590 81.640 157.350 81.920 ;
        RECT 158.470 81.640 163.790 81.920 ;
        RECT 152.870 81.360 157.350 81.640 ;
        RECT 158.750 81.360 163.790 81.640 ;
        RECT 152.870 81.080 157.630 81.360 ;
        RECT 159.030 81.080 163.790 81.360 ;
        RECT 153.150 80.800 157.910 81.080 ;
        RECT 159.310 80.800 163.790 81.080 ;
        RECT 153.430 80.520 158.190 80.800 ;
        RECT 159.590 80.520 163.790 80.800 ;
        RECT 176.950 81.640 181.430 81.920 ;
        RECT 182.550 81.640 187.310 81.920 ;
        RECT 222.310 81.640 225.950 82.200 ;
        RECT 236.310 81.920 237.990 82.760 ;
        RECT 238.550 82.760 240.510 83.040 ;
        RECT 243.870 82.760 260.390 83.040 ;
        RECT 238.550 81.920 240.790 82.760 ;
        RECT 243.870 82.480 260.670 82.760 ;
        RECT 244.150 82.200 260.950 82.480 ;
        RECT 244.150 81.920 271.590 82.200 ;
        RECT 236.310 81.640 238.270 81.920 ;
        RECT 176.950 81.360 181.150 81.640 ;
        RECT 182.550 81.360 187.030 81.640 ;
        RECT 176.950 81.080 180.870 81.360 ;
        RECT 182.270 81.080 187.030 81.360 ;
        RECT 222.030 81.080 225.670 81.640 ;
        RECT 176.950 80.800 180.590 81.080 ;
        RECT 181.990 80.800 186.750 81.080 ;
        RECT 176.950 80.520 180.310 80.800 ;
        RECT 181.710 80.520 186.470 80.800 ;
        RECT 221.750 80.520 225.390 81.080 ;
        RECT 236.590 80.800 238.270 81.640 ;
        RECT 238.830 81.640 240.790 81.920 ;
        RECT 244.430 81.640 271.590 81.920 ;
        RECT 238.830 81.080 241.070 81.640 ;
        RECT 244.430 81.360 260.110 81.640 ;
        RECT 239.110 80.800 241.070 81.080 ;
        RECT 244.710 81.080 260.110 81.360 ;
        RECT 244.710 80.800 259.830 81.080 ;
        RECT 153.710 80.240 158.470 80.520 ;
        RECT 159.870 80.240 163.790 80.520 ;
        RECT 176.670 80.240 180.030 80.520 ;
        RECT 181.430 80.240 186.190 80.520 ;
        RECT 221.470 80.240 225.110 80.520 ;
        RECT 153.710 79.960 159.030 80.240 ;
        RECT 160.150 79.960 164.070 80.240 ;
        RECT 176.110 79.960 179.750 80.240 ;
        RECT 180.870 79.960 186.190 80.240 ;
        RECT 221.190 79.960 225.110 80.240 ;
        RECT 236.870 79.960 238.550 80.800 ;
        RECT 239.110 79.960 241.350 80.800 ;
        RECT 244.990 80.520 248.630 80.800 ;
        RECT 243.310 80.240 246.670 80.520 ;
        RECT 248.350 80.240 248.630 80.520 ;
        RECT 249.470 80.240 259.550 80.800 ;
        RECT 242.470 79.960 243.870 80.240 ;
        RECT 245.830 79.960 246.390 80.240 ;
        RECT 248.350 79.960 248.910 80.240 ;
        RECT 153.990 79.680 159.310 79.960 ;
        RECT 160.710 79.680 164.350 79.960 ;
        RECT 175.550 79.680 179.190 79.960 ;
        RECT 180.590 79.680 185.910 79.960 ;
        RECT 221.190 79.680 224.830 79.960 ;
        RECT 236.870 79.680 238.830 79.960 ;
        RECT 154.270 79.400 159.590 79.680 ;
        RECT 160.990 79.400 164.910 79.680 ;
        RECT 174.990 79.400 178.910 79.680 ;
        RECT 180.310 79.400 185.630 79.680 ;
        RECT 220.910 79.400 224.830 79.680 ;
        RECT 154.550 79.120 159.870 79.400 ;
        RECT 161.550 79.120 165.750 79.400 ;
        RECT 174.150 79.120 178.350 79.400 ;
        RECT 180.030 79.120 185.350 79.400 ;
        RECT 220.910 79.120 224.550 79.400 ;
        RECT 154.830 78.840 160.430 79.120 ;
        RECT 162.110 78.840 166.870 79.120 ;
        RECT 173.030 78.840 177.790 79.120 ;
        RECT 179.470 78.840 185.070 79.120 ;
        RECT 209.150 78.840 211.670 79.120 ;
        RECT 220.630 78.840 224.550 79.120 ;
        RECT 237.150 78.840 238.830 79.680 ;
        RECT 239.390 79.680 241.350 79.960 ;
        RECT 241.630 79.680 242.750 79.960 ;
        RECT 239.390 79.400 242.190 79.680 ;
        RECT 239.390 79.120 241.630 79.400 ;
        RECT 246.110 79.120 246.670 79.960 ;
        RECT 239.390 78.840 241.350 79.120 ;
        RECT 246.390 78.840 246.670 79.120 ;
        RECT 155.110 78.560 160.710 78.840 ;
        RECT 162.390 78.560 168.550 78.840 ;
        RECT 171.350 78.560 177.510 78.840 ;
        RECT 179.190 78.560 184.790 78.840 ;
        RECT 206.630 78.560 214.190 78.840 ;
        RECT 220.630 78.560 224.270 78.840 ;
        RECT 237.150 78.560 239.110 78.840 ;
        RECT 155.390 78.280 161.270 78.560 ;
        RECT 162.950 78.280 176.950 78.560 ;
        RECT 178.630 78.280 184.510 78.560 ;
        RECT 205.230 78.280 209.430 78.560 ;
        RECT 211.390 78.280 215.870 78.560 ;
        RECT 220.350 78.280 224.270 78.560 ;
        RECT 155.670 78.000 161.830 78.280 ;
        RECT 163.790 78.000 176.110 78.280 ;
        RECT 178.070 78.000 184.230 78.280 ;
        RECT 204.390 78.000 206.910 78.280 ;
        RECT 213.910 78.000 216.990 78.280 ;
        RECT 220.350 78.000 223.990 78.280 ;
        RECT 155.950 77.720 162.110 78.000 ;
        RECT 164.350 77.720 175.550 78.000 ;
        RECT 177.790 77.720 183.950 78.000 ;
        RECT 203.550 77.720 205.790 78.000 ;
        RECT 215.310 77.720 217.830 78.000 ;
        RECT 220.070 77.720 223.990 78.000 ;
        RECT 156.230 77.440 162.670 77.720 ;
        RECT 165.190 77.440 174.710 77.720 ;
        RECT 177.230 77.440 183.670 77.720 ;
        RECT 202.710 77.440 204.670 77.720 ;
        RECT 216.430 77.440 218.670 77.720 ;
        RECT 220.070 77.440 223.710 77.720 ;
        RECT 237.430 77.440 239.110 78.560 ;
        RECT 239.670 78.560 241.070 78.840 ;
        RECT 239.670 78.280 240.790 78.560 ;
        RECT 246.110 78.280 246.670 78.840 ;
        RECT 248.630 78.280 248.910 79.960 ;
        RECT 249.470 79.960 270.750 80.240 ;
        RECT 249.470 79.680 270.470 79.960 ;
        RECT 249.190 79.120 260.110 79.400 ;
        RECT 239.670 78.000 240.510 78.280 ;
        RECT 246.110 78.000 246.390 78.280 ;
        RECT 239.670 77.440 240.230 78.000 ;
        RECT 244.990 77.720 246.390 78.000 ;
        RECT 248.350 77.720 248.910 78.280 ;
        RECT 258.990 78.000 259.550 78.280 ;
        RECT 249.190 77.720 270.750 78.000 ;
        RECT 243.870 77.440 248.630 77.720 ;
        RECT 156.510 77.160 163.510 77.440 ;
        RECT 166.310 77.160 173.590 77.440 ;
        RECT 176.390 77.160 183.390 77.440 ;
        RECT 202.150 77.160 203.830 77.440 ;
        RECT 217.550 77.160 219.510 77.440 ;
        RECT 219.790 77.160 223.430 77.440 ;
        RECT 156.790 76.880 164.070 77.160 ;
        RECT 167.990 76.880 171.910 77.160 ;
        RECT 175.830 76.880 183.110 77.160 ;
        RECT 201.590 76.880 202.990 77.160 ;
        RECT 218.390 76.880 223.430 77.160 ;
        RECT 157.070 76.600 164.910 76.880 ;
        RECT 174.990 76.600 182.830 76.880 ;
        RECT 201.310 76.600 202.430 76.880 ;
        RECT 219.230 76.600 223.150 76.880 ;
        RECT 157.630 76.320 166.030 76.600 ;
        RECT 173.870 76.320 182.270 76.600 ;
        RECT 201.310 76.320 202.150 76.600 ;
        RECT 219.510 76.320 223.150 76.600 ;
        RECT 237.710 76.600 238.830 77.440 ;
        RECT 239.670 77.160 239.950 77.440 ;
        RECT 243.310 77.160 244.990 77.440 ;
        RECT 247.510 77.160 248.630 77.440 ;
        RECT 258.990 77.440 270.750 77.720 ;
        RECT 239.390 76.880 239.950 77.160 ;
        RECT 242.750 76.880 244.150 77.160 ;
        RECT 247.230 76.880 248.070 77.160 ;
        RECT 258.990 76.880 259.550 77.440 ;
        RECT 239.390 76.600 239.670 76.880 ;
        RECT 242.470 76.600 243.590 76.880 ;
        RECT 247.230 76.600 247.790 76.880 ;
        RECT 252.830 76.600 253.390 76.880 ;
        RECT 255.350 76.600 256.190 76.880 ;
        RECT 237.710 76.320 238.550 76.600 ;
        RECT 157.910 76.040 167.150 76.320 ;
        RECT 172.750 76.040 181.990 76.320 ;
        RECT 201.590 76.040 202.990 76.320 ;
        RECT 158.190 75.760 181.710 76.040 ;
        RECT 201.870 75.760 204.390 76.040 ;
        RECT 219.230 75.760 222.870 76.320 ;
        RECT 158.750 75.480 181.150 75.760 ;
        RECT 202.430 75.480 209.990 75.760 ;
        RECT 218.950 75.480 222.870 75.760 ;
        RECT 237.990 75.480 238.550 76.320 ;
        RECT 159.310 75.200 180.590 75.480 ;
        RECT 201.870 75.200 212.230 75.480 ;
        RECT 218.950 75.200 223.430 75.480 ;
        RECT 238.270 75.200 238.550 75.480 ;
        RECT 239.110 76.040 239.670 76.600 ;
        RECT 242.190 76.320 243.030 76.600 ;
        RECT 242.190 76.040 242.750 76.320 ;
        RECT 246.950 76.040 247.510 76.600 ;
        RECT 249.750 76.320 250.590 76.600 ;
        RECT 252.830 76.320 253.670 76.600 ;
        RECT 255.350 76.320 256.470 76.600 ;
        RECT 159.590 74.920 180.310 75.200 ;
        RECT 201.310 74.920 213.910 75.200 ;
        RECT 218.670 74.920 223.710 75.200 ;
        RECT 160.150 74.640 179.750 74.920 ;
        RECT 200.750 74.640 215.030 74.920 ;
        RECT 218.670 74.640 222.310 74.920 ;
        RECT 222.870 74.640 223.990 74.920 ;
        RECT 238.270 74.640 238.550 74.920 ;
        RECT 160.710 74.360 179.190 74.640 ;
        RECT 200.190 74.360 216.150 74.640 ;
        RECT 161.270 74.080 178.630 74.360 ;
        RECT 199.630 74.080 216.990 74.360 ;
        RECT 218.390 74.080 222.030 74.640 ;
        RECT 223.430 74.360 224.550 74.640 ;
        RECT 223.710 74.080 224.830 74.360 ;
        RECT 161.830 73.800 178.070 74.080 ;
        RECT 199.070 73.800 217.830 74.080 ;
        RECT 218.110 73.800 221.750 74.080 ;
        RECT 224.270 73.800 225.110 74.080 ;
        RECT 162.670 73.520 177.230 73.800 ;
        RECT 198.790 73.520 221.750 73.800 ;
        RECT 224.550 73.520 225.390 73.800 ;
        RECT 239.110 73.520 239.390 76.040 ;
        RECT 241.910 75.760 242.750 76.040 ;
        RECT 241.910 75.200 242.470 75.760 ;
        RECT 241.910 74.080 242.750 75.200 ;
        RECT 246.670 74.080 247.230 76.040 ;
        RECT 249.750 75.760 250.870 76.320 ;
        RECT 252.830 76.040 253.950 76.320 ;
        RECT 255.350 76.040 256.750 76.320 ;
        RECT 252.830 75.760 254.230 76.040 ;
        RECT 255.630 75.760 257.030 76.040 ;
        RECT 250.030 75.480 251.150 75.760 ;
        RECT 253.110 75.480 254.230 75.760 ;
        RECT 255.910 75.480 257.030 75.760 ;
        RECT 259.270 75.480 259.830 76.880 ;
        RECT 250.030 75.200 251.430 75.480 ;
        RECT 250.310 74.920 251.430 75.200 ;
        RECT 253.390 74.920 254.510 75.480 ;
        RECT 256.190 74.920 257.030 75.480 ;
        RECT 259.550 74.920 260.110 75.480 ;
        RECT 250.590 74.640 251.430 74.920 ;
        RECT 253.950 74.640 254.230 74.920 ;
        RECT 259.550 74.640 260.950 74.920 ;
        RECT 251.150 74.360 251.430 74.640 ;
        RECT 259.550 74.360 271.310 74.640 ;
        RECT 257.590 74.080 263.750 74.360 ;
        RECT 241.910 73.800 243.030 74.080 ;
        RECT 163.510 73.240 176.390 73.520 ;
        RECT 198.230 73.240 221.470 73.520 ;
        RECT 224.830 73.240 225.670 73.520 ;
        RECT 164.350 72.960 175.550 73.240 ;
        RECT 197.950 72.960 208.310 73.240 ;
        RECT 212.230 72.960 221.470 73.240 ;
        RECT 225.110 72.960 225.950 73.240 ;
        RECT 239.110 72.960 239.670 73.520 ;
        RECT 242.190 73.240 243.030 73.800 ;
        RECT 246.950 73.240 247.510 74.080 ;
        RECT 254.790 73.800 257.030 74.080 ;
        RECT 259.830 73.800 260.390 74.080 ;
        RECT 251.990 73.520 254.230 73.800 ;
        RECT 260.110 73.520 260.670 73.800 ;
        RECT 249.190 73.240 251.430 73.520 ;
        RECT 260.110 73.240 260.950 73.520 ;
        RECT 165.470 72.680 174.430 72.960 ;
        RECT 197.390 72.680 206.630 72.960 ;
        RECT 213.910 72.680 221.190 72.960 ;
        RECT 225.390 72.680 226.230 72.960 ;
        RECT 239.390 72.680 239.670 72.960 ;
        RECT 242.470 72.680 243.310 73.240 ;
        RECT 247.230 72.960 248.630 73.240 ;
        RECT 253.950 72.960 254.510 73.240 ;
        RECT 256.470 72.960 257.310 73.240 ;
        RECT 260.390 72.960 260.950 73.240 ;
        RECT 247.230 72.680 247.790 72.960 ;
        RECT 167.150 72.400 172.750 72.680 ;
        RECT 197.110 72.400 205.510 72.680 ;
        RECT 215.030 72.400 221.190 72.680 ;
        RECT 225.670 72.400 226.510 72.680 ;
        RECT 239.390 72.400 239.950 72.680 ;
        RECT 242.750 72.400 243.590 72.680 ;
        RECT 246.950 72.400 247.790 72.680 ;
        RECT 196.830 72.120 204.670 72.400 ;
        RECT 215.870 72.120 221.190 72.400 ;
        RECT 225.950 72.120 226.790 72.400 ;
        RECT 239.670 72.120 239.950 72.400 ;
        RECT 243.030 72.120 244.430 72.400 ;
        RECT 246.110 72.120 247.790 72.400 ;
        RECT 196.550 71.840 203.830 72.120 ;
        RECT 207.190 71.840 213.070 72.120 ;
        RECT 216.710 71.840 221.750 72.120 ;
        RECT 226.230 71.840 227.070 72.120 ;
        RECT 239.670 71.840 240.230 72.120 ;
        RECT 243.590 71.840 247.790 72.120 ;
        RECT 250.870 72.400 251.710 72.960 ;
        RECT 253.670 72.680 254.790 72.960 ;
        RECT 256.470 72.680 257.590 72.960 ;
        RECT 260.670 72.680 261.230 72.960 ;
        RECT 253.670 72.400 255.070 72.680 ;
        RECT 256.470 72.400 257.870 72.680 ;
        RECT 260.670 72.400 261.510 72.680 ;
        RECT 250.870 72.120 251.990 72.400 ;
        RECT 253.950 72.120 255.070 72.400 ;
        RECT 256.750 72.120 257.870 72.400 ;
        RECT 260.950 72.120 261.510 72.400 ;
        RECT 250.870 71.840 252.270 72.120 ;
        RECT 195.990 71.560 202.990 71.840 ;
        RECT 206.070 71.560 214.470 71.840 ;
        RECT 216.990 71.560 222.310 71.840 ;
        RECT 226.510 71.560 227.350 71.840 ;
        RECT 239.950 71.560 240.510 71.840 ;
        RECT 244.430 71.560 245.830 71.840 ;
        RECT 195.710 71.280 202.430 71.560 ;
        RECT 204.950 71.280 215.310 71.560 ;
        RECT 216.710 71.280 222.590 71.560 ;
        RECT 195.430 71.000 201.870 71.280 ;
        RECT 204.110 71.000 216.150 71.280 ;
        RECT 216.710 71.000 222.870 71.280 ;
        RECT 226.790 71.000 227.630 71.560 ;
        RECT 239.950 71.280 240.790 71.560 ;
        RECT 247.230 71.280 247.790 71.840 ;
        RECT 251.150 71.560 252.550 71.840 ;
        RECT 254.230 71.560 255.350 72.120 ;
        RECT 257.030 71.560 258.150 72.120 ;
        RECT 261.230 71.840 261.790 72.120 ;
        RECT 261.230 71.560 262.070 71.840 ;
        RECT 251.430 71.280 252.550 71.560 ;
        RECT 254.510 71.280 255.350 71.560 ;
        RECT 257.310 71.280 258.150 71.560 ;
        RECT 261.510 71.280 262.070 71.560 ;
        RECT 240.230 71.000 241.070 71.280 ;
        RECT 247.230 71.000 248.070 71.280 ;
        RECT 251.710 71.000 252.550 71.280 ;
        RECT 255.070 71.000 255.350 71.280 ;
        RECT 261.790 71.000 262.350 71.280 ;
        RECT 195.150 70.720 201.590 71.000 ;
        RECT 203.550 70.720 223.430 71.000 ;
        RECT 227.070 70.720 227.910 71.000 ;
        RECT 239.110 70.720 239.390 71.000 ;
        RECT 240.510 70.720 241.350 71.000 ;
        RECT 194.870 70.440 201.030 70.720 ;
        RECT 202.990 70.440 223.710 70.720 ;
        RECT 227.350 70.440 228.190 70.720 ;
        RECT 194.590 70.160 200.470 70.440 ;
        RECT 202.430 70.160 208.310 70.440 ;
        RECT 194.310 69.880 200.190 70.160 ;
        RECT 201.870 69.880 207.470 70.160 ;
        RECT 210.270 69.880 210.830 70.440 ;
        RECT 212.230 70.160 223.990 70.440 ;
        RECT 227.630 70.160 228.190 70.440 ;
        RECT 239.110 70.440 239.670 70.720 ;
        RECT 241.070 70.440 241.630 70.720 ;
        RECT 247.510 70.440 248.070 71.000 ;
        RECT 261.790 70.720 262.630 71.000 ;
        RECT 261.510 70.440 262.630 70.720 ;
        RECT 239.110 70.160 239.950 70.440 ;
        RECT 241.350 70.160 242.190 70.440 ;
        RECT 247.510 70.160 248.350 70.440 ;
        RECT 257.590 70.160 262.910 70.440 ;
        RECT 123.470 69.600 131.310 69.880 ;
        RECT 135.790 69.600 138.590 69.880 ;
        RECT 140.550 69.600 143.350 69.880 ;
        RECT 146.150 69.600 148.950 69.880 ;
        RECT 151.190 69.600 153.990 69.880 ;
        RECT 156.510 69.600 159.590 69.880 ;
        RECT 194.030 69.600 199.910 69.880 ;
        RECT 201.310 69.600 205.790 69.880 ;
        RECT 126.830 69.320 135.510 69.600 ;
        RECT 128.790 68.480 135.510 69.320 ;
        RECT 128.510 67.920 135.230 68.480 ;
        RECT 137.190 68.200 139.150 69.600 ;
        RECT 137.190 67.920 138.870 68.200 ;
        RECT 141.950 67.920 145.030 69.600 ;
        RECT 147.550 69.320 150.630 69.600 ;
        RECT 148.670 68.760 150.630 69.320 ;
        RECT 148.670 68.480 150.350 68.760 ;
        RECT 130.750 66.800 132.710 67.920 ;
        RECT 136.910 66.800 138.870 67.920 ;
        RECT 130.750 66.520 132.430 66.800 ;
        RECT 136.910 66.520 138.590 66.800 ;
        RECT 141.670 66.520 145.030 67.920 ;
        RECT 148.390 67.360 150.350 68.480 ;
        RECT 152.310 67.920 154.270 69.600 ;
        RECT 157.910 69.320 160.430 69.600 ;
        RECT 194.030 69.320 199.350 69.600 ;
        RECT 201.030 69.320 204.950 69.600 ;
        RECT 158.470 69.040 160.430 69.320 ;
        RECT 193.750 69.040 199.070 69.320 ;
        RECT 200.470 69.040 204.670 69.320 ;
        RECT 158.190 68.480 160.150 69.040 ;
        RECT 193.470 68.760 198.790 69.040 ;
        RECT 200.190 68.760 203.830 69.040 ;
        RECT 204.390 68.760 204.670 69.040 ;
        RECT 193.190 68.480 198.510 68.760 ;
        RECT 199.910 68.480 203.270 68.760 ;
        RECT 157.910 67.920 159.870 68.480 ;
        RECT 192.910 68.200 198.230 68.480 ;
        RECT 199.350 68.200 202.710 68.480 ;
        RECT 202.990 68.200 203.550 68.480 ;
        RECT 204.390 68.200 204.950 68.760 ;
        RECT 192.910 67.920 197.950 68.200 ;
        RECT 199.070 67.920 202.150 68.200 ;
        RECT 203.270 67.920 203.830 68.200 ;
        RECT 152.590 67.360 154.270 67.920 ;
        RECT 157.630 67.360 159.590 67.920 ;
        RECT 192.630 67.640 197.670 67.920 ;
        RECT 198.790 67.640 201.870 67.920 ;
        RECT 203.550 67.640 204.390 67.920 ;
        RECT 204.670 67.640 204.950 68.200 ;
        RECT 192.350 67.360 197.390 67.640 ;
        RECT 198.510 67.360 201.310 67.640 ;
        RECT 203.830 67.360 204.950 67.640 ;
        RECT 148.390 67.080 150.070 67.360 ;
        RECT 130.470 65.400 132.430 66.520 ;
        RECT 136.630 65.400 138.590 66.520 ;
        RECT 141.390 66.240 145.030 66.520 ;
        RECT 141.390 65.960 143.350 66.240 ;
        RECT 141.390 65.400 143.070 65.960 ;
        RECT 130.470 65.120 132.150 65.400 ;
        RECT 130.190 64.000 132.150 65.120 ;
        RECT 136.350 64.280 138.310 65.400 ;
        RECT 141.110 64.280 143.070 65.400 ;
        RECT 136.350 64.000 138.030 64.280 ;
        RECT 141.110 64.000 142.790 64.280 ;
        RECT 130.190 63.720 131.870 64.000 ;
        RECT 129.910 62.880 131.870 63.720 ;
        RECT 136.070 62.880 138.030 64.000 ;
        RECT 140.830 62.880 142.790 64.000 ;
        RECT 143.630 62.880 145.030 66.240 ;
        RECT 148.110 65.960 150.070 67.080 ;
        RECT 147.830 64.840 149.790 65.960 ;
        RECT 147.830 64.560 149.510 64.840 ;
        RECT 147.550 63.440 149.510 64.560 ;
        RECT 152.590 64.280 154.550 67.360 ;
        RECT 157.630 67.080 159.310 67.360 ;
        RECT 192.350 67.080 197.110 67.360 ;
        RECT 198.230 67.080 201.030 67.360 ;
        RECT 204.390 67.080 205.230 67.360 ;
        RECT 157.350 66.800 159.310 67.080 ;
        RECT 192.070 66.800 196.830 67.080 ;
        RECT 197.950 66.800 201.590 67.080 ;
        RECT 204.670 66.800 205.230 67.080 ;
        RECT 157.350 66.520 159.030 66.800 ;
        RECT 157.070 66.240 159.030 66.520 ;
        RECT 191.790 66.520 196.550 66.800 ;
        RECT 197.670 66.520 200.470 66.800 ;
        RECT 201.030 66.520 201.870 66.800 ;
        RECT 204.670 66.520 205.510 66.800 ;
        RECT 191.790 66.240 196.270 66.520 ;
        RECT 197.390 66.240 200.190 66.520 ;
        RECT 201.590 66.240 202.430 66.520 ;
        RECT 204.950 66.240 206.070 66.520 ;
        RECT 157.070 65.960 158.750 66.240 ;
        RECT 156.790 65.680 158.750 65.960 ;
        RECT 191.510 65.680 195.990 66.240 ;
        RECT 197.390 65.960 199.910 66.240 ;
        RECT 201.870 65.960 202.710 66.240 ;
        RECT 197.110 65.680 199.630 65.960 ;
        RECT 202.430 65.680 203.270 65.960 ;
        RECT 204.950 65.680 205.230 66.240 ;
        RECT 205.510 65.960 206.350 66.240 ;
        RECT 206.910 65.960 207.190 69.880 ;
        RECT 210.550 69.320 210.830 69.880 ;
        RECT 212.790 69.880 213.350 70.160 ;
        RECT 213.630 69.880 219.790 70.160 ;
        RECT 220.350 69.880 224.270 70.160 ;
        RECT 227.630 69.880 228.470 70.160 ;
        RECT 239.390 69.880 240.510 70.160 ;
        RECT 241.630 69.880 242.750 70.160 ;
        RECT 247.230 69.880 248.630 70.160 ;
        RECT 253.670 69.880 260.950 70.160 ;
        RECT 212.790 69.600 213.070 69.880 ;
        RECT 213.910 69.600 214.470 69.880 ;
        RECT 214.750 69.600 219.790 69.880 ;
        RECT 220.630 69.600 224.830 69.880 ;
        RECT 227.910 69.600 228.750 69.880 ;
        RECT 210.550 68.760 211.110 69.320 ;
        RECT 212.790 69.040 213.350 69.600 ;
        RECT 213.630 69.320 214.190 69.600 ;
        RECT 215.310 69.320 219.510 69.600 ;
        RECT 220.910 69.320 225.110 69.600 ;
        RECT 228.190 69.320 228.750 69.600 ;
        RECT 239.390 69.600 240.790 69.880 ;
        RECT 241.910 69.600 243.310 69.880 ;
        RECT 246.390 69.600 247.510 69.880 ;
        RECT 248.070 69.600 248.910 69.880 ;
        RECT 249.750 69.600 258.990 69.880 ;
        RECT 239.390 69.320 241.350 69.600 ;
        RECT 241.910 69.320 246.950 69.600 ;
        RECT 248.350 69.320 259.270 69.600 ;
        RECT 213.630 69.040 213.910 69.320 ;
        RECT 212.790 68.760 213.910 69.040 ;
        RECT 215.590 69.040 219.790 69.320 ;
        RECT 221.470 69.040 225.390 69.320 ;
        RECT 228.190 69.040 229.030 69.320 ;
        RECT 215.590 68.760 220.350 69.040 ;
        RECT 221.750 68.760 225.670 69.040 ;
        RECT 228.470 68.760 229.030 69.040 ;
        RECT 210.830 68.200 211.110 68.760 ;
        RECT 213.070 68.200 213.630 68.760 ;
        RECT 215.310 68.480 220.630 68.760 ;
        RECT 222.030 68.480 225.950 68.760 ;
        RECT 228.470 68.480 229.310 68.760 ;
        RECT 215.310 68.200 220.910 68.480 ;
        RECT 222.310 68.200 225.950 68.480 ;
        RECT 228.750 68.200 229.310 68.480 ;
        RECT 239.670 68.200 241.630 69.320 ;
        RECT 241.910 69.040 245.550 69.320 ;
        RECT 248.630 69.040 254.510 69.320 ;
        RECT 255.070 69.040 259.830 69.320 ;
        RECT 242.190 68.760 244.150 69.040 ;
        RECT 248.350 68.760 250.310 69.040 ;
        RECT 250.590 68.760 254.230 69.040 ;
        RECT 255.350 68.760 258.710 69.040 ;
        RECT 259.270 68.760 260.390 69.040 ;
        RECT 210.830 67.360 211.390 68.200 ;
        RECT 212.790 67.920 213.350 68.200 ;
        RECT 212.510 67.360 213.350 67.920 ;
        RECT 215.030 67.920 221.190 68.200 ;
        RECT 222.590 67.920 226.230 68.200 ;
        RECT 228.750 67.920 229.590 68.200 ;
        RECT 215.030 67.640 221.470 67.920 ;
        RECT 222.870 67.640 226.510 67.920 ;
        RECT 229.030 67.640 229.590 67.920 ;
        RECT 211.110 66.800 211.390 67.360 ;
        RECT 212.230 67.080 212.790 67.360 ;
        RECT 211.110 66.520 211.670 66.800 ;
        RECT 211.950 66.520 212.510 67.080 ;
        RECT 211.110 66.240 212.230 66.520 ;
        RECT 213.070 66.240 213.630 67.360 ;
        RECT 214.750 67.080 218.670 67.640 ;
        RECT 218.950 67.360 221.750 67.640 ;
        RECT 223.150 67.360 226.790 67.640 ;
        RECT 229.030 67.360 229.870 67.640 ;
        RECT 239.950 67.360 241.910 68.200 ;
        RECT 242.190 67.920 244.430 68.760 ;
        RECT 248.070 68.200 250.030 68.760 ;
        RECT 250.870 68.480 254.510 68.760 ;
        RECT 255.070 68.480 258.430 68.760 ;
        RECT 259.270 68.480 260.670 68.760 ;
        RECT 250.870 68.200 258.710 68.480 ;
        RECT 259.270 68.200 260.950 68.480 ;
        RECT 247.790 67.920 250.310 68.200 ;
        RECT 250.590 67.920 261.230 68.200 ;
        RECT 219.230 67.080 222.030 67.360 ;
        RECT 223.430 67.080 227.070 67.360 ;
        RECT 214.470 66.800 218.390 67.080 ;
        RECT 219.790 66.800 222.310 67.080 ;
        RECT 223.710 66.800 227.070 67.080 ;
        RECT 229.310 67.080 229.870 67.360 ;
        RECT 240.230 67.080 241.910 67.360 ;
        RECT 242.470 67.640 244.430 67.920 ;
        RECT 247.510 67.640 261.790 67.920 ;
        RECT 242.470 67.080 244.710 67.640 ;
        RECT 247.230 67.360 250.030 67.640 ;
        RECT 251.150 67.360 262.070 67.640 ;
        RECT 229.310 66.800 230.150 67.080 ;
        RECT 214.190 66.520 218.390 66.800 ;
        RECT 220.070 66.520 222.590 66.800 ;
        RECT 223.990 66.520 227.350 66.800 ;
        RECT 229.590 66.520 230.150 66.800 ;
        RECT 240.230 66.520 242.190 67.080 ;
        RECT 214.190 66.240 218.110 66.520 ;
        RECT 208.590 65.960 213.630 66.240 ;
        RECT 213.910 65.960 218.110 66.240 ;
        RECT 220.070 66.240 222.870 66.520 ;
        RECT 223.990 66.240 227.630 66.520 ;
        RECT 229.590 66.240 230.430 66.520 ;
        RECT 220.070 65.960 223.150 66.240 ;
        RECT 224.270 65.960 227.910 66.240 ;
        RECT 206.070 65.680 206.630 65.960 ;
        RECT 206.910 65.680 217.830 65.960 ;
        RECT 156.790 65.400 158.470 65.680 ;
        RECT 156.510 65.120 158.470 65.400 ;
        RECT 191.230 65.400 195.710 65.680 ;
        RECT 196.830 65.400 199.350 65.680 ;
        RECT 202.710 65.400 203.550 65.680 ;
        RECT 191.230 65.120 195.430 65.400 ;
        RECT 156.510 64.840 158.190 65.120 ;
        RECT 156.230 64.560 158.190 64.840 ;
        RECT 190.950 64.840 195.430 65.120 ;
        RECT 196.550 65.120 199.070 65.400 ;
        RECT 203.270 65.120 204.110 65.400 ;
        RECT 204.950 65.120 205.510 65.680 ;
        RECT 206.350 65.400 217.830 65.680 ;
        RECT 219.790 65.400 220.350 65.960 ;
        RECT 220.910 65.680 223.430 65.960 ;
        RECT 224.550 65.680 227.910 65.960 ;
        RECT 229.870 65.680 230.430 66.240 ;
        RECT 240.510 65.960 242.190 66.520 ;
        RECT 242.750 66.800 244.710 67.080 ;
        RECT 246.950 67.080 249.190 67.360 ;
        RECT 251.710 67.080 262.350 67.360 ;
        RECT 246.950 66.800 248.910 67.080 ;
        RECT 250.030 66.800 250.870 67.080 ;
        RECT 251.990 66.800 262.350 67.080 ;
        RECT 242.750 65.960 244.990 66.800 ;
        RECT 221.190 65.400 223.710 65.680 ;
        RECT 206.350 65.120 217.550 65.400 ;
        RECT 219.510 65.120 223.710 65.400 ;
        RECT 224.830 65.120 228.190 65.680 ;
        RECT 229.870 65.400 230.710 65.680 ;
        RECT 240.510 65.400 242.470 65.960 ;
        RECT 196.550 64.840 198.790 65.120 ;
        RECT 203.550 64.840 204.390 65.120 ;
        RECT 205.230 64.840 205.510 65.120 ;
        RECT 205.790 64.840 209.150 65.120 ;
        RECT 212.790 64.840 217.550 65.120 ;
        RECT 219.230 64.840 220.910 65.120 ;
        RECT 221.750 64.840 223.990 65.120 ;
        RECT 225.110 64.840 228.470 65.120 ;
        RECT 230.150 64.840 230.710 65.400 ;
        RECT 190.950 64.560 195.150 64.840 ;
        RECT 196.270 64.560 198.510 64.840 ;
        RECT 204.110 64.560 204.950 64.840 ;
        RECT 205.230 64.560 208.030 64.840 ;
        RECT 213.350 64.560 217.270 64.840 ;
        RECT 218.670 64.560 220.070 64.840 ;
        RECT 221.750 64.560 224.270 64.840 ;
        RECT 225.110 64.560 228.750 64.840 ;
        RECT 230.150 64.560 230.990 64.840 ;
        RECT 240.790 64.560 242.470 65.400 ;
        RECT 243.030 65.680 244.990 65.960 ;
        RECT 246.670 66.520 247.230 66.800 ;
        RECT 247.510 66.520 248.630 66.800 ;
        RECT 249.470 66.520 251.430 66.800 ;
        RECT 252.270 66.520 261.510 66.800 ;
        RECT 261.790 66.520 262.630 66.800 ;
        RECT 246.670 65.960 246.950 66.520 ;
        RECT 247.790 66.240 248.630 66.520 ;
        RECT 249.190 66.240 251.710 66.520 ;
        RECT 247.790 65.960 248.350 66.240 ;
        RECT 246.670 65.680 248.350 65.960 ;
        RECT 243.030 64.840 245.270 65.680 ;
        RECT 246.950 64.840 248.350 65.680 ;
        RECT 243.310 64.560 245.270 64.840 ;
        RECT 156.230 64.280 157.910 64.560 ;
        RECT 147.550 63.160 149.230 63.440 ;
        RECT 129.910 62.600 131.590 62.880 ;
        RECT 136.070 62.600 137.750 62.880 ;
        RECT 140.830 62.600 142.510 62.880 ;
        RECT 129.630 61.480 131.590 62.600 ;
        RECT 135.790 61.480 137.750 62.600 ;
        RECT 140.550 61.480 142.510 62.600 ;
        RECT 129.630 61.200 131.310 61.480 ;
        RECT 135.790 61.200 137.470 61.480 ;
        RECT 140.550 61.200 142.230 61.480 ;
        RECT 129.350 60.080 131.310 61.200 ;
        RECT 135.510 60.360 137.470 61.200 ;
        RECT 140.270 60.360 142.230 61.200 ;
        RECT 135.510 60.080 137.190 60.360 ;
        RECT 140.270 60.080 141.950 60.360 ;
        RECT 129.350 59.800 131.030 60.080 ;
        RECT 129.070 58.680 131.030 59.800 ;
        RECT 135.230 58.960 137.190 60.080 ;
        RECT 139.990 58.960 141.950 60.080 ;
        RECT 143.630 59.520 145.310 62.880 ;
        RECT 147.270 62.040 149.230 63.160 ;
        RECT 146.990 60.920 148.950 62.040 ;
        RECT 152.870 61.480 154.550 64.280 ;
        RECT 155.950 64.000 157.910 64.280 ;
        RECT 190.670 64.280 195.150 64.560 ;
        RECT 195.990 64.280 198.510 64.560 ;
        RECT 204.390 64.280 207.190 64.560 ;
        RECT 213.070 64.280 217.270 64.560 ;
        RECT 217.830 64.280 219.510 64.560 ;
        RECT 222.030 64.280 224.270 64.560 ;
        RECT 225.390 64.280 228.750 64.560 ;
        RECT 190.670 64.000 194.870 64.280 ;
        RECT 195.990 64.000 198.790 64.280 ;
        RECT 204.390 64.000 206.630 64.280 ;
        RECT 213.070 64.000 218.390 64.280 ;
        RECT 218.950 64.000 219.230 64.280 ;
        RECT 222.310 64.000 224.550 64.280 ;
        RECT 155.950 63.720 157.630 64.000 ;
        RECT 155.670 63.440 157.630 63.720 ;
        RECT 190.390 63.440 194.590 64.000 ;
        RECT 195.710 63.720 197.950 64.000 ;
        RECT 198.510 63.720 199.070 64.000 ;
        RECT 204.110 63.720 206.070 64.000 ;
        RECT 195.710 63.440 197.670 63.720 ;
        RECT 198.790 63.440 199.350 63.720 ;
        RECT 203.830 63.440 205.790 63.720 ;
        RECT 212.790 63.440 217.830 64.000 ;
        RECT 218.670 63.720 219.230 64.000 ;
        RECT 222.590 63.720 224.550 64.000 ;
        RECT 225.670 63.720 229.030 64.280 ;
        RECT 230.430 63.720 230.990 64.560 ;
        RECT 218.670 63.440 218.950 63.720 ;
        RECT 155.670 63.160 157.350 63.440 ;
        RECT 190.390 63.160 194.310 63.440 ;
        RECT 155.390 62.880 157.350 63.160 ;
        RECT 190.110 62.880 194.310 63.160 ;
        RECT 195.430 63.160 197.670 63.440 ;
        RECT 195.430 62.880 197.390 63.160 ;
        RECT 199.070 62.880 199.630 63.440 ;
        RECT 203.550 63.160 205.230 63.440 ;
        RECT 212.510 63.160 218.110 63.440 ;
        RECT 218.390 63.160 218.950 63.440 ;
        RECT 222.590 63.160 224.830 63.720 ;
        RECT 225.950 63.160 229.310 63.720 ;
        RECT 230.430 63.440 231.270 63.720 ;
        RECT 241.070 63.440 242.750 64.560 ;
        RECT 243.310 63.720 245.550 64.560 ;
        RECT 247.230 64.280 248.350 64.840 ;
        RECT 248.910 64.560 251.990 66.240 ;
        RECT 252.550 65.960 261.230 66.520 ;
        RECT 262.070 65.960 262.630 66.520 ;
        RECT 252.550 65.680 262.630 65.960 ;
        RECT 252.550 64.560 262.350 65.680 ;
        RECT 249.190 64.280 251.710 64.560 ;
        RECT 252.550 64.280 254.230 64.560 ;
        RECT 258.150 64.280 262.350 64.560 ;
        RECT 247.510 64.000 248.630 64.280 ;
        RECT 249.470 64.000 251.710 64.280 ;
        RECT 252.270 64.000 254.230 64.280 ;
        RECT 254.790 64.000 257.870 64.280 ;
        RECT 247.510 63.720 248.910 64.000 ;
        RECT 249.750 63.720 251.150 64.000 ;
        RECT 252.270 63.720 254.510 64.000 ;
        RECT 254.790 63.720 257.590 64.000 ;
        RECT 258.150 63.720 262.070 64.280 ;
        RECT 243.590 63.440 245.550 63.720 ;
        RECT 247.790 63.440 249.190 63.720 ;
        RECT 251.710 63.440 254.510 63.720 ;
        RECT 203.270 62.880 204.950 63.160 ;
        RECT 212.510 62.880 218.670 63.160 ;
        RECT 221.190 62.880 225.110 63.160 ;
        RECT 155.390 62.320 157.070 62.880 ;
        RECT 190.110 62.600 194.030 62.880 ;
        RECT 155.110 61.760 156.790 62.320 ;
        RECT 189.830 62.040 194.030 62.600 ;
        RECT 195.150 62.600 197.390 62.880 ;
        RECT 199.350 62.600 199.910 62.880 ;
        RECT 202.990 62.600 204.670 62.880 ;
        RECT 209.990 62.600 211.670 62.880 ;
        RECT 212.230 62.600 218.670 62.880 ;
        RECT 219.510 62.600 222.030 62.880 ;
        RECT 223.150 62.600 225.110 62.880 ;
        RECT 226.230 62.600 229.590 63.160 ;
        RECT 230.710 62.600 231.270 63.440 ;
        RECT 241.350 62.600 243.030 63.440 ;
        RECT 243.590 62.600 245.830 63.440 ;
        RECT 247.790 63.160 249.470 63.440 ;
        RECT 251.430 63.160 254.790 63.440 ;
        RECT 255.070 63.160 257.310 63.720 ;
        RECT 257.870 63.440 262.070 63.720 ;
        RECT 257.870 63.160 261.790 63.440 ;
        RECT 248.070 62.880 254.790 63.160 ;
        RECT 255.350 62.880 257.030 63.160 ;
        RECT 257.590 62.880 260.390 63.160 ;
        RECT 260.950 62.880 261.790 63.160 ;
        RECT 195.150 62.320 197.110 62.600 ;
        RECT 199.630 62.320 200.190 62.600 ;
        RECT 202.710 62.320 204.390 62.600 ;
        RECT 208.590 62.320 221.470 62.600 ;
        RECT 194.870 62.040 197.110 62.320 ;
        RECT 199.910 62.040 200.470 62.320 ;
        RECT 202.430 62.040 204.110 62.320 ;
        RECT 208.030 62.040 221.470 62.320 ;
        RECT 223.430 62.040 225.390 62.600 ;
        RECT 226.510 62.320 229.870 62.600 ;
        RECT 230.710 62.320 231.550 62.600 ;
        RECT 226.510 62.040 230.150 62.320 ;
        RECT 152.870 61.200 154.270 61.480 ;
        RECT 155.110 61.200 156.510 61.760 ;
        RECT 189.830 61.480 193.750 62.040 ;
        RECT 194.870 61.760 197.390 62.040 ;
        RECT 200.190 61.760 200.750 62.040 ;
        RECT 202.430 61.760 203.830 62.040 ;
        RECT 207.470 61.760 210.270 62.040 ;
        RECT 211.390 61.760 221.750 62.040 ;
        RECT 194.590 61.480 197.670 61.760 ;
        RECT 200.190 61.480 201.030 61.760 ;
        RECT 152.870 60.920 156.230 61.200 ;
        RECT 146.990 60.640 148.670 60.920 ;
        RECT 152.870 60.640 155.950 60.920 ;
        RECT 135.230 58.680 136.910 58.960 ;
        RECT 139.990 58.680 141.670 58.960 ;
        RECT 128.790 57.560 130.750 58.680 ;
        RECT 134.950 57.560 136.910 58.680 ;
        RECT 139.710 57.560 141.670 58.680 ;
        RECT 128.790 57.280 130.470 57.560 ;
        RECT 134.950 57.280 136.630 57.560 ;
        RECT 139.710 57.280 141.390 57.560 ;
        RECT 128.510 56.160 130.470 57.280 ;
        RECT 134.670 56.440 136.630 57.280 ;
        RECT 139.430 56.440 141.390 57.280 ;
        RECT 134.670 56.160 136.350 56.440 ;
        RECT 139.430 56.160 141.110 56.440 ;
        RECT 128.510 55.880 130.190 56.160 ;
        RECT 128.230 54.760 130.190 55.880 ;
        RECT 134.390 55.040 136.350 56.160 ;
        RECT 139.150 55.040 141.110 56.160 ;
        RECT 134.390 54.760 136.070 55.040 ;
        RECT 139.150 54.760 140.830 55.040 ;
        RECT 128.230 54.480 129.910 54.760 ;
        RECT 127.950 53.640 129.910 54.480 ;
        RECT 134.110 53.640 136.070 54.760 ;
        RECT 138.870 53.640 140.830 54.760 ;
        RECT 143.910 54.760 145.310 59.520 ;
        RECT 146.710 59.520 148.670 60.640 ;
        RECT 153.150 60.360 155.950 60.640 ;
        RECT 189.550 60.640 193.470 61.480 ;
        RECT 194.590 60.920 196.550 61.480 ;
        RECT 197.390 61.200 197.950 61.480 ;
        RECT 200.470 61.200 201.030 61.480 ;
        RECT 202.150 61.200 203.550 61.760 ;
        RECT 206.910 61.480 209.150 61.760 ;
        RECT 211.670 61.480 215.590 61.760 ;
        RECT 216.150 61.480 221.750 61.760 ;
        RECT 206.630 61.200 208.310 61.480 ;
        RECT 211.670 61.200 215.310 61.480 ;
        RECT 216.710 61.200 221.750 61.480 ;
        RECT 223.710 61.480 225.670 62.040 ;
        RECT 226.510 61.760 230.430 62.040 ;
        RECT 226.790 61.480 230.710 61.760 ;
        RECT 230.990 61.480 231.550 62.320 ;
        RECT 241.630 61.480 243.310 62.600 ;
        RECT 243.870 62.320 245.830 62.600 ;
        RECT 248.350 62.600 255.070 62.880 ;
        RECT 248.350 62.320 249.190 62.600 ;
        RECT 249.750 62.320 255.070 62.600 ;
        RECT 255.630 62.600 257.030 62.880 ;
        RECT 257.310 62.600 260.110 62.880 ;
        RECT 255.630 62.320 256.750 62.600 ;
        RECT 257.310 62.320 260.390 62.600 ;
        RECT 260.950 62.320 261.510 62.880 ;
        RECT 243.870 61.480 246.110 62.320 ;
        RECT 248.630 62.040 248.910 62.320 ;
        RECT 249.750 62.040 255.350 62.320 ;
        RECT 255.910 62.040 256.750 62.320 ;
        RECT 257.030 62.040 261.510 62.320 ;
        RECT 248.630 61.760 249.190 62.040 ;
        RECT 249.750 61.760 255.630 62.040 ;
        RECT 255.910 61.760 256.470 62.040 ;
        RECT 257.030 61.760 261.230 62.040 ;
        RECT 248.910 61.480 255.630 61.760 ;
        RECT 256.750 61.480 261.230 61.760 ;
        RECT 223.710 61.200 225.950 61.480 ;
        RECT 197.670 60.920 198.230 61.200 ;
        RECT 200.750 60.920 201.310 61.200 ;
        RECT 201.870 60.920 203.270 61.200 ;
        RECT 206.350 60.920 207.750 61.200 ;
        RECT 211.390 60.920 215.310 61.200 ;
        RECT 189.550 60.360 193.190 60.640 ;
        RECT 153.150 59.800 155.670 60.360 ;
        RECT 146.710 59.240 148.390 59.520 ;
        RECT 146.430 58.120 148.390 59.240 ;
        RECT 153.150 59.240 155.390 59.800 ;
        RECT 189.270 59.520 193.190 60.360 ;
        RECT 194.310 60.360 196.270 60.920 ;
        RECT 197.950 60.640 198.510 60.920 ;
        RECT 201.030 60.640 202.990 60.920 ;
        RECT 206.070 60.640 207.470 60.920 ;
        RECT 211.390 60.640 215.590 60.920 ;
        RECT 216.990 60.640 221.470 61.200 ;
        RECT 223.990 60.920 225.950 61.200 ;
        RECT 226.790 60.920 231.550 61.480 ;
        RECT 223.710 60.640 225.950 60.920 ;
        RECT 227.070 60.640 231.550 60.920 ;
        RECT 241.910 61.200 243.310 61.480 ;
        RECT 244.150 61.200 246.110 61.480 ;
        RECT 249.190 61.200 255.910 61.480 ;
        RECT 256.470 61.200 260.950 61.480 ;
        RECT 241.910 60.640 243.590 61.200 ;
        RECT 198.230 60.360 199.070 60.640 ;
        RECT 201.310 60.360 202.990 60.640 ;
        RECT 205.790 60.360 207.190 60.640 ;
        RECT 211.110 60.360 215.870 60.640 ;
        RECT 216.710 60.360 221.190 60.640 ;
        RECT 223.150 60.360 226.230 60.640 ;
        RECT 194.310 60.080 202.710 60.360 ;
        RECT 205.510 60.080 206.630 60.360 ;
        RECT 209.430 60.080 216.150 60.360 ;
        RECT 216.430 60.080 221.470 60.360 ;
        RECT 222.870 60.080 223.710 60.360 ;
        RECT 194.030 59.800 196.270 60.080 ;
        RECT 198.790 59.800 199.910 60.080 ;
        RECT 200.750 59.800 202.710 60.080 ;
        RECT 153.150 58.400 155.110 59.240 ;
        RECT 189.270 58.960 192.910 59.520 ;
        RECT 153.150 58.120 154.830 58.400 ;
        RECT 146.150 57.000 148.110 58.120 ;
        RECT 152.870 57.000 154.830 58.120 ;
        RECT 188.990 57.840 192.910 58.960 ;
        RECT 194.030 59.240 195.990 59.800 ;
        RECT 199.350 59.520 199.910 59.800 ;
        RECT 201.310 59.520 202.430 59.800 ;
        RECT 205.230 59.520 206.350 60.080 ;
        RECT 208.870 59.800 209.710 60.080 ;
        RECT 210.830 59.800 214.750 60.080 ;
        RECT 215.310 59.800 221.470 60.080 ;
        RECT 222.310 59.800 223.150 60.080 ;
        RECT 208.310 59.660 209.010 59.800 ;
        RECT 208.310 59.520 208.870 59.660 ;
        RECT 199.630 59.240 200.190 59.520 ;
        RECT 201.030 59.240 202.430 59.520 ;
        RECT 204.950 59.240 206.070 59.520 ;
        RECT 208.030 59.240 208.590 59.520 ;
        RECT 194.030 58.680 195.710 59.240 ;
        RECT 199.910 58.960 200.470 59.240 ;
        RECT 201.030 58.960 202.150 59.240 ;
        RECT 200.190 58.680 202.150 58.960 ;
        RECT 193.750 57.840 195.710 58.680 ;
        RECT 200.470 58.400 202.150 58.680 ;
        RECT 204.670 58.680 205.790 59.240 ;
        RECT 207.750 58.960 208.590 59.240 ;
        RECT 210.830 59.240 214.470 59.800 ;
        RECT 215.590 59.520 222.590 59.800 ;
        RECT 224.270 59.520 226.230 60.360 ;
        RECT 227.070 60.360 231.830 60.640 ;
        RECT 227.070 60.080 230.990 60.360 ;
        RECT 227.350 59.800 230.990 60.080 ;
        RECT 242.190 60.080 243.590 60.640 ;
        RECT 244.150 60.360 246.390 61.200 ;
        RECT 249.190 60.920 260.950 61.200 ;
        RECT 249.470 60.640 260.670 60.920 ;
        RECT 249.470 60.360 260.390 60.640 ;
        RECT 244.430 60.080 246.390 60.360 ;
        RECT 249.750 60.080 260.390 60.360 ;
        RECT 242.190 59.800 243.870 60.080 ;
        RECT 215.590 59.240 222.310 59.520 ;
        RECT 224.270 59.240 226.510 59.520 ;
        RECT 210.830 58.960 214.750 59.240 ;
        RECT 215.590 58.960 222.590 59.240 ;
        RECT 207.470 58.680 208.870 58.960 ;
        RECT 211.110 58.680 222.870 58.960 ;
        RECT 204.670 58.400 205.510 58.680 ;
        RECT 207.190 58.400 207.750 58.680 ;
        RECT 208.310 58.400 209.150 58.680 ;
        RECT 199.630 58.120 201.870 58.400 ;
        RECT 196.830 57.840 201.870 58.120 ;
        RECT 146.150 56.720 147.830 57.000 ;
        RECT 152.870 56.720 154.550 57.000 ;
        RECT 145.870 55.600 147.830 56.720 ;
        RECT 152.590 55.600 154.550 56.720 ;
        RECT 145.870 55.040 147.550 55.600 ;
        RECT 152.590 55.320 154.270 55.600 ;
        RECT 145.590 54.760 147.550 55.040 ;
        RECT 143.910 54.200 147.550 54.760 ;
        RECT 152.310 54.200 154.270 55.320 ;
        RECT 127.950 53.360 129.630 53.640 ;
        RECT 134.110 53.360 135.790 53.640 ;
        RECT 138.870 53.360 140.550 53.640 ;
        RECT 127.670 52.240 129.630 53.360 ;
        RECT 133.830 52.240 135.790 53.360 ;
        RECT 138.590 52.240 140.550 53.360 ;
        RECT 143.910 52.800 147.270 54.200 ;
        RECT 152.030 53.080 153.990 54.200 ;
        RECT 188.990 53.360 192.630 57.840 ;
        RECT 193.750 57.560 197.950 57.840 ;
        RECT 193.750 57.280 195.710 57.560 ;
        RECT 193.750 54.480 195.430 57.280 ;
        RECT 200.750 57.000 201.870 57.840 ;
        RECT 204.390 58.120 205.510 58.400 ;
        RECT 206.910 58.120 207.470 58.400 ;
        RECT 208.590 58.120 209.430 58.400 ;
        RECT 211.390 58.120 222.870 58.680 ;
        RECT 224.550 58.400 226.510 59.240 ;
        RECT 227.350 58.960 231.270 59.800 ;
        RECT 242.470 58.960 243.870 59.800 ;
        RECT 244.430 59.520 246.670 60.080 ;
        RECT 250.030 59.800 260.110 60.080 ;
        RECT 244.710 59.240 246.670 59.520 ;
        RECT 250.310 59.520 258.150 59.800 ;
        RECT 258.710 59.520 259.830 59.800 ;
        RECT 250.310 59.240 251.710 59.520 ;
        RECT 251.990 59.240 257.870 59.520 ;
        RECT 258.990 59.240 259.550 59.520 ;
        RECT 224.270 58.120 226.510 58.400 ;
        RECT 204.390 57.560 205.230 58.120 ;
        RECT 206.910 57.840 207.190 58.120 ;
        RECT 208.870 57.840 209.710 58.120 ;
        RECT 200.470 56.720 201.870 57.000 ;
        RECT 204.110 57.280 205.230 57.560 ;
        RECT 206.630 57.560 207.190 57.840 ;
        RECT 209.150 57.560 209.990 57.840 ;
        RECT 211.390 57.560 211.950 58.120 ;
        RECT 212.230 57.840 213.350 58.120 ;
        RECT 213.910 57.840 222.870 58.120 ;
        RECT 223.710 57.840 226.510 58.120 ;
        RECT 227.630 57.840 231.270 58.960 ;
        RECT 242.750 58.400 244.150 58.960 ;
        RECT 244.710 58.400 246.950 59.240 ;
        RECT 250.590 58.960 251.430 59.240 ;
        RECT 250.870 58.680 251.430 58.960 ;
        RECT 252.270 58.960 258.150 59.240 ;
        RECT 258.710 58.960 259.550 59.240 ;
        RECT 252.270 58.680 259.270 58.960 ;
        RECT 251.150 58.400 258.990 58.680 ;
        RECT 243.030 57.840 244.150 58.400 ;
        RECT 244.990 58.120 246.950 58.400 ;
        RECT 251.430 58.120 258.710 58.400 ;
        RECT 214.470 57.560 222.590 57.840 ;
        RECT 223.150 57.560 223.990 57.840 ;
        RECT 200.470 55.320 201.590 56.720 ;
        RECT 200.470 55.040 201.870 55.320 ;
        RECT 193.750 54.200 196.830 54.480 ;
        RECT 193.750 53.920 198.230 54.200 ;
        RECT 200.750 53.920 201.870 55.040 ;
        RECT 204.110 54.760 204.950 57.280 ;
        RECT 206.630 56.720 206.910 57.560 ;
        RECT 209.430 57.280 211.950 57.560 ;
        RECT 209.710 57.000 211.950 57.280 ;
        RECT 209.710 56.720 210.550 57.000 ;
        RECT 211.110 56.720 211.950 57.000 ;
        RECT 214.750 57.280 223.430 57.560 ;
        RECT 214.750 56.720 222.870 57.280 ;
        RECT 224.830 56.720 226.790 57.840 ;
        RECT 227.630 56.720 231.550 57.840 ;
        RECT 243.030 57.560 244.430 57.840 ;
        RECT 243.310 56.720 244.430 57.560 ;
        RECT 244.990 57.560 247.230 58.120 ;
        RECT 247.510 57.840 248.910 58.120 ;
        RECT 251.710 57.840 258.430 58.120 ;
        RECT 247.510 57.560 247.790 57.840 ;
        RECT 248.770 57.700 249.470 57.840 ;
        RECT 248.910 57.560 249.470 57.700 ;
        RECT 251.990 57.560 257.870 57.840 ;
        RECT 244.990 57.420 247.650 57.560 ;
        RECT 249.330 57.420 250.310 57.560 ;
        RECT 244.990 57.280 247.510 57.420 ;
        RECT 249.470 57.280 250.310 57.420 ;
        RECT 252.270 57.280 257.590 57.560 ;
        RECT 206.350 56.440 206.910 56.720 ;
        RECT 206.350 55.600 206.630 56.440 ;
        RECT 209.430 55.600 209.990 56.720 ;
        RECT 211.670 56.440 212.230 56.720 ;
        RECT 211.670 56.160 212.510 56.440 ;
        RECT 214.750 56.160 222.030 56.720 ;
        RECT 222.310 56.440 223.990 56.720 ;
        RECT 225.110 56.440 226.790 56.720 ;
        RECT 223.430 56.160 226.790 56.440 ;
        RECT 211.670 55.880 214.190 56.160 ;
        RECT 214.750 55.880 222.310 56.160 ;
        RECT 224.550 55.880 226.790 56.160 ;
        RECT 211.670 55.600 222.590 55.880 ;
        RECT 206.350 55.320 206.910 55.600 ;
        RECT 209.430 55.320 210.270 55.600 ;
        RECT 211.670 55.320 212.230 55.600 ;
        RECT 214.470 55.320 222.590 55.600 ;
        RECT 204.110 54.480 205.230 54.760 ;
        RECT 204.390 53.920 205.230 54.480 ;
        RECT 206.630 54.480 206.910 55.320 ;
        RECT 209.150 55.040 210.550 55.320 ;
        RECT 211.110 55.040 211.950 55.320 ;
        RECT 208.590 54.760 211.950 55.040 ;
        RECT 214.750 55.040 215.310 55.320 ;
        RECT 215.590 55.040 222.590 55.320 ;
        RECT 208.310 54.480 209.430 54.760 ;
        RECT 210.550 54.480 211.670 54.760 ;
        RECT 214.750 54.480 215.030 55.040 ;
        RECT 215.870 54.760 222.590 55.040 ;
        RECT 206.630 54.200 207.190 54.480 ;
        RECT 207.750 54.200 208.870 54.480 ;
        RECT 206.910 53.920 208.310 54.200 ;
        RECT 152.030 52.800 153.710 53.080 ;
        RECT 127.670 51.960 129.350 52.240 ;
        RECT 127.390 51.400 129.350 51.960 ;
        RECT 133.550 51.400 135.510 52.240 ;
        RECT 138.310 51.400 140.270 52.240 ;
        RECT 143.910 51.680 146.990 52.800 ;
        RECT 151.750 51.680 153.710 52.800 ;
        RECT 188.990 52.240 192.910 53.360 ;
        RECT 193.750 52.800 195.710 53.920 ;
        RECT 196.830 53.640 199.630 53.920 ;
        RECT 200.750 53.640 202.150 53.920 ;
        RECT 204.390 53.640 205.510 53.920 ;
        RECT 206.910 53.640 207.750 53.920 ;
        RECT 198.230 53.360 202.150 53.640 ;
        RECT 199.630 53.080 202.150 53.360 ;
        RECT 204.670 53.360 205.510 53.640 ;
        RECT 207.190 53.360 207.750 53.640 ;
        RECT 204.670 53.080 205.790 53.360 ;
        RECT 207.470 53.080 208.030 53.360 ;
        RECT 211.390 53.080 211.950 54.480 ;
        RECT 214.470 54.200 215.030 54.480 ;
        RECT 216.430 54.480 222.590 54.760 ;
        RECT 225.110 54.480 226.790 55.880 ;
        RECT 227.910 54.480 231.550 56.720 ;
        RECT 243.590 56.160 244.710 56.720 ;
        RECT 245.270 56.160 247.510 57.280 ;
        RECT 250.030 57.000 250.870 57.280 ;
        RECT 252.550 57.000 254.230 57.280 ;
        RECT 250.730 56.860 251.430 57.000 ;
        RECT 250.870 56.720 251.430 56.860 ;
        RECT 252.830 56.720 254.230 57.000 ;
        RECT 255.070 57.000 257.310 57.280 ;
        RECT 255.070 56.720 256.750 57.000 ;
        RECT 251.290 56.580 251.990 56.720 ;
        RECT 251.430 56.440 251.990 56.580 ;
        RECT 253.390 56.440 256.190 56.720 ;
        RECT 251.850 56.300 252.550 56.440 ;
        RECT 251.990 56.160 252.550 56.300 ;
        RECT 253.670 56.160 255.630 56.440 ;
        RECT 243.870 55.600 244.710 56.160 ;
        RECT 245.550 55.880 247.510 56.160 ;
        RECT 252.410 56.020 253.390 56.160 ;
        RECT 252.550 55.880 253.390 56.020 ;
        RECT 254.230 55.880 255.070 56.160 ;
        RECT 243.870 55.320 244.990 55.600 ;
        RECT 244.150 54.760 244.990 55.320 ;
        RECT 245.550 55.040 247.790 55.880 ;
        RECT 253.250 55.740 254.370 55.880 ;
        RECT 253.250 55.600 254.230 55.740 ;
        RECT 250.030 55.320 250.310 55.600 ;
        RECT 251.710 55.320 251.990 55.600 ;
        RECT 253.110 55.320 253.390 55.600 ;
        RECT 254.090 55.460 255.630 55.600 ;
        RECT 254.230 55.320 255.630 55.460 ;
        RECT 245.830 54.760 248.070 55.040 ;
        RECT 249.750 54.760 250.590 55.320 ;
        RECT 251.430 55.040 252.270 55.320 ;
        RECT 251.430 54.760 251.990 55.040 ;
        RECT 252.830 54.760 253.670 55.320 ;
        RECT 255.350 55.040 258.150 55.320 ;
        RECT 258.010 54.900 258.710 55.040 ;
        RECT 258.150 54.760 258.710 54.900 ;
        RECT 244.150 54.480 245.270 54.760 ;
        RECT 245.830 54.480 248.350 54.760 ;
        RECT 258.570 54.620 258.990 54.760 ;
        RECT 258.710 54.480 258.990 54.620 ;
        RECT 216.430 54.200 222.870 54.480 ;
        RECT 214.470 53.920 214.750 54.200 ;
        RECT 216.430 53.920 217.270 54.200 ;
        RECT 217.830 53.920 221.750 54.200 ;
        RECT 222.310 53.920 223.430 54.200 ;
        RECT 214.190 53.640 214.750 53.920 ;
        RECT 213.910 53.360 214.470 53.640 ;
        RECT 216.150 53.360 217.270 53.920 ;
        RECT 219.790 53.640 220.910 53.920 ;
        RECT 223.150 53.640 223.990 53.920 ;
        RECT 213.630 53.080 214.190 53.360 ;
        RECT 200.750 52.800 202.150 53.080 ;
        RECT 204.950 52.800 205.790 53.080 ;
        RECT 207.750 52.800 208.310 53.080 ;
        RECT 193.750 52.520 195.990 52.800 ;
        RECT 200.750 52.520 202.430 52.800 ;
        RECT 204.950 52.520 206.070 52.800 ;
        RECT 208.030 52.520 208.590 52.800 ;
        RECT 189.270 51.960 192.910 52.240 ;
        RECT 143.910 51.400 146.710 51.680 ;
        RECT 151.750 51.400 153.430 51.680 ;
        RECT 189.270 50.840 193.190 51.960 ;
        RECT 194.030 51.680 195.990 52.520 ;
        RECT 200.470 52.240 202.430 52.520 ;
        RECT 205.230 52.240 206.350 52.520 ;
        RECT 208.310 52.240 209.150 52.520 ;
        RECT 211.670 52.240 212.230 53.080 ;
        RECT 213.350 52.800 213.910 53.080 ;
        RECT 215.870 52.800 216.990 53.360 ;
        RECT 219.510 53.080 220.910 53.640 ;
        RECT 223.710 53.360 224.550 53.640 ;
        RECT 224.830 53.360 226.790 54.480 ;
        RECT 227.630 53.360 231.550 54.480 ;
        RECT 244.430 53.920 245.270 54.480 ;
        RECT 246.110 54.200 248.630 54.480 ;
        RECT 246.110 53.920 248.910 54.200 ;
        RECT 250.590 53.920 251.430 54.480 ;
        RECT 252.270 53.920 253.110 54.480 ;
        RECT 253.950 54.200 254.510 54.480 ;
        RECT 258.850 54.340 259.270 54.480 ;
        RECT 258.990 54.200 259.270 54.340 ;
        RECT 253.670 53.920 254.510 54.200 ;
        RECT 259.130 54.060 259.550 54.200 ;
        RECT 259.270 53.920 259.550 54.060 ;
        RECT 244.430 53.640 245.550 53.920 ;
        RECT 244.710 53.360 245.550 53.640 ;
        RECT 246.390 53.640 249.470 53.920 ;
        RECT 250.870 53.640 251.150 53.920 ;
        RECT 252.550 53.640 252.830 53.920 ;
        RECT 253.950 53.640 254.230 53.920 ;
        RECT 259.270 53.640 259.830 53.920 ;
        RECT 246.390 53.360 250.310 53.640 ;
        RECT 259.270 53.360 260.110 53.640 ;
        RECT 224.270 53.080 226.510 53.360 ;
        RECT 219.510 52.800 220.630 53.080 ;
        RECT 213.070 52.520 213.630 52.800 ;
        RECT 215.590 52.520 216.710 52.800 ;
        RECT 212.510 52.240 213.350 52.520 ;
        RECT 200.190 51.960 202.710 52.240 ;
        RECT 205.230 51.960 206.630 52.240 ;
        RECT 208.870 51.960 209.710 52.240 ;
        RECT 211.670 51.960 212.790 52.240 ;
        RECT 215.310 51.960 216.430 52.520 ;
        RECT 219.230 52.240 220.630 52.800 ;
        RECT 224.830 52.520 226.510 53.080 ;
        RECT 227.630 52.520 231.270 53.360 ;
        RECT 244.990 53.080 245.550 53.360 ;
        RECT 246.670 53.080 265.710 53.360 ;
        RECT 244.990 52.800 245.830 53.080 ;
        RECT 246.950 52.800 265.710 53.080 ;
        RECT 245.270 52.520 246.110 52.800 ;
        RECT 247.230 52.520 265.710 52.800 ;
        RECT 199.630 51.680 202.710 51.960 ;
        RECT 205.510 51.680 206.910 51.960 ;
        RECT 209.430 51.680 212.230 51.960 ;
        RECT 215.030 51.680 216.150 51.960 ;
        RECT 218.950 51.680 220.350 52.240 ;
        RECT 224.550 51.680 226.510 52.520 ;
        RECT 194.030 51.400 196.270 51.680 ;
        RECT 196.550 51.400 202.990 51.680 ;
        RECT 205.790 51.400 207.190 51.680 ;
        RECT 214.750 51.400 215.870 51.680 ;
        RECT 218.670 51.400 220.070 51.680 ;
        RECT 224.550 51.400 226.230 51.680 ;
        RECT 194.310 51.120 200.190 51.400 ;
        RECT 201.590 51.120 202.990 51.400 ;
        RECT 206.070 51.120 207.470 51.400 ;
        RECT 214.190 51.120 215.590 51.400 ;
        RECT 218.670 51.120 222.030 51.400 ;
        RECT 224.270 51.120 226.230 51.400 ;
        RECT 227.350 51.400 231.270 52.520 ;
        RECT 245.550 52.240 246.390 52.520 ;
        RECT 247.510 52.240 265.710 52.520 ;
        RECT 245.550 51.960 246.670 52.240 ;
        RECT 248.070 51.960 265.710 52.240 ;
        RECT 245.830 51.680 246.950 51.960 ;
        RECT 248.630 51.680 265.710 51.960 ;
        RECT 246.110 51.400 247.230 51.680 ;
        RECT 249.470 51.400 265.710 51.680 ;
        RECT 227.350 51.120 230.990 51.400 ;
        RECT 246.390 51.120 247.790 51.400 ;
        RECT 189.550 50.000 193.470 50.840 ;
        RECT 194.310 50.280 196.270 51.120 ;
        RECT 199.070 50.840 199.910 51.120 ;
        RECT 201.870 50.840 203.270 51.120 ;
        RECT 206.350 50.840 207.750 51.120 ;
        RECT 213.910 50.840 215.310 51.120 ;
        RECT 218.390 50.840 220.070 51.120 ;
        RECT 221.190 50.840 226.230 51.120 ;
        RECT 198.790 50.560 199.630 50.840 ;
        RECT 201.870 50.560 203.550 50.840 ;
        RECT 206.630 50.560 208.310 50.840 ;
        RECT 213.350 50.560 215.030 50.840 ;
        RECT 218.110 50.560 220.070 50.840 ;
        RECT 198.510 50.280 199.350 50.560 ;
        RECT 201.590 50.280 203.550 50.560 ;
        RECT 206.910 50.280 209.150 50.560 ;
        RECT 212.510 50.280 214.750 50.560 ;
        RECT 218.110 50.280 219.510 50.560 ;
        RECT 219.790 50.280 220.350 50.560 ;
        RECT 189.550 49.720 193.750 50.000 ;
        RECT 189.830 49.160 193.750 49.720 ;
        RECT 194.590 49.720 196.550 50.280 ;
        RECT 198.230 50.000 199.070 50.280 ;
        RECT 201.310 50.000 202.150 50.280 ;
        RECT 202.430 50.000 203.830 50.280 ;
        RECT 207.470 50.000 210.550 50.280 ;
        RECT 211.110 50.000 214.190 50.280 ;
        RECT 217.830 50.000 219.230 50.280 ;
        RECT 220.070 50.000 220.630 50.280 ;
        RECT 223.990 50.000 225.950 50.840 ;
        RECT 227.070 50.280 230.990 51.120 ;
        RECT 246.950 50.840 248.630 51.120 ;
        RECT 247.230 50.560 249.750 50.840 ;
        RECT 247.790 50.280 263.470 50.560 ;
        RECT 197.950 49.720 198.790 50.000 ;
        RECT 201.030 49.720 201.870 50.000 ;
        RECT 202.710 49.720 204.110 50.000 ;
        RECT 208.030 49.720 213.630 50.000 ;
        RECT 217.550 49.720 219.230 50.000 ;
        RECT 194.590 49.440 196.830 49.720 ;
        RECT 197.670 49.440 198.510 49.720 ;
        RECT 200.750 49.440 201.590 49.720 ;
        RECT 202.710 49.440 204.390 49.720 ;
        RECT 208.870 49.440 213.070 49.720 ;
        RECT 217.270 49.440 219.510 49.720 ;
        RECT 220.350 49.440 220.910 50.000 ;
        RECT 223.710 49.440 225.670 50.000 ;
        RECT 226.790 49.440 230.710 50.280 ;
        RECT 248.630 50.000 263.470 50.280 ;
        RECT 194.870 49.160 196.830 49.440 ;
        RECT 197.390 49.160 198.230 49.440 ;
        RECT 200.470 49.160 201.310 49.440 ;
        RECT 202.990 49.160 204.670 49.440 ;
        RECT 210.270 49.160 211.390 49.440 ;
        RECT 216.990 49.160 221.190 49.440 ;
        RECT 223.430 49.160 225.670 49.440 ;
        RECT 226.510 49.160 230.710 49.440 ;
        RECT 189.830 48.880 194.030 49.160 ;
        RECT 194.870 48.880 197.950 49.160 ;
        RECT 200.190 48.880 201.030 49.160 ;
        RECT 203.270 48.880 204.950 49.160 ;
        RECT 216.710 48.880 218.950 49.160 ;
        RECT 220.070 48.880 222.310 49.160 ;
        RECT 223.430 48.880 225.390 49.160 ;
        RECT 226.510 48.880 230.430 49.160 ;
        RECT 190.110 48.600 194.030 48.880 ;
        RECT 195.150 48.600 197.670 48.880 ;
        RECT 200.190 48.600 200.750 48.880 ;
        RECT 203.550 48.600 205.510 48.880 ;
        RECT 216.430 48.600 218.110 48.880 ;
        RECT 138.310 48.320 145.870 48.600 ;
        RECT 157.350 48.320 159.870 48.600 ;
        RECT 166.590 48.320 169.110 48.600 ;
        RECT 174.990 48.320 177.510 48.600 ;
        RECT 181.150 48.320 183.390 48.600 ;
        RECT 139.430 48.040 148.670 48.320 ;
        RECT 150.910 48.040 152.590 48.320 ;
        RECT 157.910 48.040 163.230 48.320 ;
        RECT 166.870 48.040 173.030 48.320 ;
        RECT 175.270 48.040 178.910 48.320 ;
        RECT 181.710 48.040 184.790 48.320 ;
        RECT 190.110 48.040 194.310 48.600 ;
        RECT 195.150 48.320 197.390 48.600 ;
        RECT 199.910 48.320 200.470 48.600 ;
        RECT 203.830 48.320 205.790 48.600 ;
        RECT 215.870 48.320 217.830 48.600 ;
        RECT 218.670 48.320 219.230 48.880 ;
        RECT 221.190 48.600 225.390 48.880 ;
        RECT 221.470 48.320 222.030 48.600 ;
        RECT 142.790 47.200 148.670 48.040 ;
        RECT 142.790 46.640 148.390 47.200 ;
        RECT 150.630 46.920 152.590 48.040 ;
        RECT 159.590 47.760 163.230 48.040 ;
        RECT 168.550 47.760 173.310 48.040 ;
        RECT 159.870 47.480 163.230 47.760 ;
        RECT 168.270 47.480 173.310 47.760 ;
        RECT 150.630 46.640 152.310 46.920 ;
        RECT 159.590 46.640 163.230 47.480 ;
        RECT 167.990 47.200 173.590 47.480 ;
        RECT 167.710 46.920 173.870 47.200 ;
        RECT 176.950 46.920 178.910 48.040 ;
        RECT 182.830 47.760 184.790 48.040 ;
        RECT 190.390 47.760 194.310 48.040 ;
        RECT 195.430 48.040 197.390 48.320 ;
        RECT 199.630 48.040 200.470 48.320 ;
        RECT 204.110 48.040 206.350 48.320 ;
        RECT 215.590 48.040 217.550 48.320 ;
        RECT 218.950 48.040 219.510 48.320 ;
        RECT 221.470 48.040 222.310 48.320 ;
        RECT 195.430 47.760 197.670 48.040 ;
        RECT 199.350 47.760 200.190 48.040 ;
        RECT 204.390 47.760 206.630 48.040 ;
        RECT 215.030 47.760 217.270 48.040 ;
        RECT 219.230 47.760 219.510 48.040 ;
        RECT 221.750 47.760 222.310 48.040 ;
        RECT 222.870 48.040 225.110 48.600 ;
        RECT 226.230 48.320 230.430 48.880 ;
        RECT 226.230 48.040 230.150 48.320 ;
        RECT 222.870 47.760 224.830 48.040 ;
        RECT 182.830 47.480 184.510 47.760 ;
        RECT 167.150 46.640 174.150 46.920 ;
        RECT 176.950 46.640 178.630 46.920 ;
        RECT 142.510 45.520 144.470 46.640 ;
        RECT 150.350 45.520 152.310 46.640 ;
        RECT 159.310 46.080 160.990 46.640 ;
        RECT 161.270 46.360 163.230 46.640 ;
        RECT 159.310 45.800 160.710 46.080 ;
        RECT 161.550 45.800 163.230 46.360 ;
        RECT 166.870 46.360 169.670 46.640 ;
        RECT 171.630 46.360 174.430 46.640 ;
        RECT 166.870 46.080 169.390 46.360 ;
        RECT 171.910 46.080 174.430 46.360 ;
        RECT 166.870 45.800 169.110 46.080 ;
        RECT 171.910 45.800 174.150 46.080 ;
        RECT 142.510 45.240 144.190 45.520 ;
        RECT 150.350 45.240 152.030 45.520 ;
        RECT 159.030 45.240 160.710 45.800 ;
        RECT 142.230 44.120 144.190 45.240 ;
        RECT 150.070 44.120 152.030 45.240 ;
        RECT 158.750 44.960 160.710 45.240 ;
        RECT 158.750 44.400 160.430 44.960 ;
        RECT 158.470 44.120 160.430 44.400 ;
        RECT 141.950 43.000 143.910 44.120 ;
        RECT 149.790 43.000 151.750 44.120 ;
        RECT 158.470 43.560 160.150 44.120 ;
        RECT 158.190 43.280 160.150 43.560 ;
        RECT 161.270 43.280 162.950 45.800 ;
        RECT 166.590 44.960 168.550 45.800 ;
        RECT 166.590 44.680 168.270 44.960 ;
        RECT 166.310 43.560 168.270 44.680 ;
        RECT 172.190 44.680 174.150 45.800 ;
        RECT 176.670 45.520 178.630 46.640 ;
        RECT 182.550 46.360 184.510 47.480 ;
        RECT 190.390 47.480 194.590 47.760 ;
        RECT 195.710 47.480 197.670 47.760 ;
        RECT 199.070 47.480 199.910 47.760 ;
        RECT 204.950 47.480 207.470 47.760 ;
        RECT 214.190 47.480 216.710 47.760 ;
        RECT 219.230 47.480 219.790 47.760 ;
        RECT 222.030 47.480 224.830 47.760 ;
        RECT 225.950 47.480 230.150 48.040 ;
        RECT 190.390 47.200 194.870 47.480 ;
        RECT 195.710 47.200 197.950 47.480 ;
        RECT 198.790 47.200 199.630 47.480 ;
        RECT 205.230 47.200 208.030 47.480 ;
        RECT 213.630 47.200 216.430 47.480 ;
        RECT 219.510 47.200 219.790 47.480 ;
        RECT 190.670 46.920 194.870 47.200 ;
        RECT 195.990 46.920 198.230 47.200 ;
        RECT 198.510 46.920 199.350 47.200 ;
        RECT 204.950 46.920 209.150 47.200 ;
        RECT 212.510 46.920 215.870 47.200 ;
        RECT 219.510 46.920 220.070 47.200 ;
        RECT 222.310 46.920 224.550 47.480 ;
        RECT 225.670 47.200 229.870 47.480 ;
        RECT 225.390 46.920 229.870 47.200 ;
        RECT 190.670 46.640 195.150 46.920 ;
        RECT 195.990 46.640 199.070 46.920 ;
        RECT 204.390 46.640 205.510 46.920 ;
        RECT 205.790 46.640 215.310 46.920 ;
        RECT 190.950 46.360 195.150 46.640 ;
        RECT 196.270 46.360 198.790 46.640 ;
        RECT 203.830 46.360 204.950 46.640 ;
        RECT 182.550 46.080 184.230 46.360 ;
        RECT 190.950 46.080 195.430 46.360 ;
        RECT 196.550 46.080 198.790 46.360 ;
        RECT 203.270 46.080 204.390 46.360 ;
        RECT 205.790 46.080 206.350 46.640 ;
        RECT 206.910 46.360 215.310 46.640 ;
        RECT 219.790 46.360 220.350 46.920 ;
        RECT 222.030 46.640 224.270 46.920 ;
        RECT 225.390 46.640 229.590 46.920 ;
        RECT 221.750 46.360 223.990 46.640 ;
        RECT 206.630 46.080 213.910 46.360 ;
        RECT 214.190 46.080 215.590 46.360 ;
        RECT 220.070 46.080 220.630 46.360 ;
        RECT 176.670 45.240 178.350 45.520 ;
        RECT 172.190 44.400 173.870 44.680 ;
        RECT 166.310 43.280 167.990 43.560 ;
        RECT 141.950 42.720 143.630 43.000 ;
        RECT 149.790 42.720 151.470 43.000 ;
        RECT 158.190 42.720 159.870 43.280 ;
        RECT 141.670 41.600 143.630 42.720 ;
        RECT 149.510 41.600 151.470 42.720 ;
        RECT 157.910 42.440 159.870 42.720 ;
        RECT 157.910 42.160 159.590 42.440 ;
        RECT 157.630 41.600 159.590 42.160 ;
        RECT 141.670 41.320 143.350 41.600 ;
        RECT 149.510 41.320 151.190 41.600 ;
        RECT 157.630 41.320 159.310 41.600 ;
        RECT 141.390 40.200 143.350 41.320 ;
        RECT 149.230 40.200 151.190 41.320 ;
        RECT 157.350 41.040 159.310 41.320 ;
        RECT 160.990 41.040 162.950 43.280 ;
        RECT 166.030 42.160 167.990 43.280 ;
        RECT 171.910 43.280 173.870 44.400 ;
        RECT 176.390 44.120 178.350 45.240 ;
        RECT 182.270 44.960 184.230 46.080 ;
        RECT 191.230 45.520 195.710 46.080 ;
        RECT 196.550 45.800 199.070 46.080 ;
        RECT 202.990 45.800 204.110 46.080 ;
        RECT 205.790 45.800 207.190 46.080 ;
        RECT 196.830 45.520 199.350 45.800 ;
        RECT 202.430 45.520 203.550 45.800 ;
        RECT 205.790 45.520 206.910 45.800 ;
        RECT 191.510 45.240 195.990 45.520 ;
        RECT 197.110 45.240 199.630 45.520 ;
        RECT 201.870 45.240 202.990 45.520 ;
        RECT 205.790 45.240 206.630 45.520 ;
        RECT 191.510 44.960 196.270 45.240 ;
        RECT 197.390 44.960 199.910 45.240 ;
        RECT 201.310 44.960 202.430 45.240 ;
        RECT 205.510 44.960 206.350 45.240 ;
        RECT 182.270 44.680 183.950 44.960 ;
        RECT 191.790 44.680 196.270 44.960 ;
        RECT 197.670 44.680 200.190 44.960 ;
        RECT 200.750 44.680 201.870 44.960 ;
        RECT 204.950 44.680 206.350 44.960 ;
        RECT 207.470 44.680 208.030 46.080 ;
        RECT 208.870 45.800 213.350 46.080 ;
        RECT 212.230 45.520 213.630 45.800 ;
        RECT 171.910 43.000 173.590 43.280 ;
        RECT 171.630 42.720 173.590 43.000 ;
        RECT 176.110 43.000 178.070 44.120 ;
        RECT 181.990 43.840 183.950 44.680 ;
        RECT 192.070 44.400 196.550 44.680 ;
        RECT 197.670 44.400 201.590 44.680 ;
        RECT 204.670 44.400 206.350 44.680 ;
        RECT 192.070 44.120 196.830 44.400 ;
        RECT 197.950 44.120 201.030 44.400 ;
        RECT 204.390 44.120 205.230 44.400 ;
        RECT 192.350 43.840 197.110 44.120 ;
        RECT 198.230 43.840 201.030 44.120 ;
        RECT 204.110 43.840 204.950 44.120 ;
        RECT 205.790 43.840 206.070 44.400 ;
        RECT 181.990 43.280 183.670 43.840 ;
        RECT 192.350 43.560 197.390 43.840 ;
        RECT 198.510 43.560 201.590 43.840 ;
        RECT 203.830 43.560 204.670 43.840 ;
        RECT 192.630 43.280 197.670 43.560 ;
        RECT 198.790 43.280 201.870 43.560 ;
        RECT 203.550 43.280 204.390 43.560 ;
        RECT 176.110 42.720 177.790 43.000 ;
        RECT 166.030 41.880 168.270 42.160 ;
        RECT 165.750 41.600 168.550 41.880 ;
        RECT 175.830 41.600 177.790 42.720 ;
        RECT 181.710 42.440 183.670 43.280 ;
        RECT 192.910 43.000 197.950 43.280 ;
        RECT 199.350 43.000 202.430 43.280 ;
        RECT 203.270 43.000 204.110 43.280 ;
        RECT 193.190 42.720 198.230 43.000 ;
        RECT 199.630 42.720 203.830 43.000 ;
        RECT 193.190 42.440 198.510 42.720 ;
        RECT 199.910 42.440 203.550 42.720 ;
        RECT 181.710 42.160 183.390 42.440 ;
        RECT 193.470 42.160 198.790 42.440 ;
        RECT 200.190 42.160 203.830 42.440 ;
        RECT 165.750 41.320 168.830 41.600 ;
        RECT 175.830 41.320 177.510 41.600 ;
        RECT 166.030 41.040 169.110 41.320 ;
        RECT 157.350 40.480 159.030 41.040 ;
        RECT 157.070 40.200 159.030 40.480 ;
        RECT 141.390 39.920 146.710 40.200 ;
        RECT 149.230 39.920 150.910 40.200 ;
        RECT 141.110 39.640 146.710 39.920 ;
        RECT 141.110 38.800 146.430 39.640 ;
        RECT 148.950 39.080 150.910 39.920 ;
        RECT 157.070 39.640 158.750 40.200 ;
        RECT 156.790 39.360 158.750 39.640 ;
        RECT 160.990 39.360 162.670 41.040 ;
        RECT 166.310 40.760 169.390 41.040 ;
        RECT 166.590 40.480 169.670 40.760 ;
        RECT 166.870 40.200 169.950 40.480 ;
        RECT 175.550 40.200 177.510 41.320 ;
        RECT 181.430 41.040 183.390 42.160 ;
        RECT 193.750 41.880 199.070 42.160 ;
        RECT 200.750 41.880 204.390 42.160 ;
        RECT 194.030 41.600 199.350 41.880 ;
        RECT 201.030 41.600 205.230 41.880 ;
        RECT 205.510 41.600 206.070 43.840 ;
        RECT 194.310 41.320 199.910 41.600 ;
        RECT 201.590 41.320 206.070 41.600 ;
        RECT 207.750 43.560 208.030 44.680 ;
        RECT 211.950 45.240 212.790 45.520 ;
        RECT 213.070 45.240 213.910 45.520 ;
        RECT 211.950 44.400 212.510 45.240 ;
        RECT 213.350 44.960 213.910 45.240 ;
        RECT 214.190 44.960 214.750 46.080 ;
        RECT 215.030 45.800 215.870 46.080 ;
        RECT 220.350 45.800 220.630 46.080 ;
        RECT 221.470 46.080 223.990 46.360 ;
        RECT 225.110 46.360 229.590 46.640 ;
        RECT 225.110 46.080 229.310 46.360 ;
        RECT 221.470 45.800 223.710 46.080 ;
        RECT 224.830 45.800 229.310 46.080 ;
        RECT 215.310 45.520 216.150 45.800 ;
        RECT 220.350 45.520 220.910 45.800 ;
        RECT 221.190 45.520 223.430 45.800 ;
        RECT 215.590 45.240 216.430 45.520 ;
        RECT 220.630 45.240 223.430 45.520 ;
        RECT 224.550 45.240 229.030 45.800 ;
        RECT 215.870 44.960 216.710 45.240 ;
        RECT 220.630 44.960 223.150 45.240 ;
        RECT 224.270 44.960 228.750 45.240 ;
        RECT 213.350 44.680 214.750 44.960 ;
        RECT 216.150 44.680 216.710 44.960 ;
        RECT 220.350 44.680 222.870 44.960 ;
        RECT 223.990 44.680 228.750 44.960 ;
        RECT 213.630 44.400 214.470 44.680 ;
        RECT 216.150 44.400 216.990 44.680 ;
        RECT 220.070 44.400 222.590 44.680 ;
        RECT 223.710 44.400 228.470 44.680 ;
        RECT 211.670 43.560 212.230 44.400 ;
        RECT 194.590 41.040 200.190 41.320 ;
        RECT 201.870 41.040 206.910 41.320 ;
        RECT 207.750 41.040 208.310 43.560 ;
        RECT 211.390 43.280 212.230 43.560 ;
        RECT 213.910 44.120 214.470 44.400 ;
        RECT 216.430 44.120 217.270 44.400 ;
        RECT 219.510 44.120 222.310 44.400 ;
        RECT 223.710 44.120 228.190 44.400 ;
        RECT 213.910 43.560 214.750 44.120 ;
        RECT 216.710 43.840 217.550 44.120 ;
        RECT 219.230 43.840 222.030 44.120 ;
        RECT 223.430 43.840 228.190 44.120 ;
        RECT 216.990 43.560 217.830 43.840 ;
        RECT 218.950 43.560 221.750 43.840 ;
        RECT 223.150 43.560 227.910 43.840 ;
        RECT 213.910 43.280 215.030 43.560 ;
        RECT 217.270 43.280 217.830 43.560 ;
        RECT 218.390 43.280 221.470 43.560 ;
        RECT 222.870 43.280 227.630 43.560 ;
        RECT 211.390 42.440 211.950 43.280 ;
        RECT 213.910 43.000 215.310 43.280 ;
        RECT 213.910 42.440 214.470 43.000 ;
        RECT 214.750 42.720 215.310 43.000 ;
        RECT 217.550 43.000 221.190 43.280 ;
        RECT 222.590 43.000 227.630 43.280 ;
        RECT 217.550 42.720 220.910 43.000 ;
        RECT 222.310 42.720 227.350 43.000 ;
        RECT 215.030 42.440 215.590 42.720 ;
        RECT 217.270 42.440 220.630 42.720 ;
        RECT 222.030 42.440 227.070 42.720 ;
        RECT 211.110 41.600 211.670 42.440 ;
        RECT 213.910 42.160 214.190 42.440 ;
        RECT 215.030 42.160 215.870 42.440 ;
        RECT 216.710 42.160 220.070 42.440 ;
        RECT 221.750 42.160 226.790 42.440 ;
        RECT 181.430 40.760 183.110 41.040 ;
        RECT 194.590 40.760 200.750 41.040 ;
        RECT 202.430 40.760 208.590 41.040 ;
        RECT 210.830 40.760 211.390 41.600 ;
        RECT 213.630 41.320 214.190 42.160 ;
        RECT 215.310 41.880 219.790 42.160 ;
        RECT 221.190 41.880 226.790 42.160 ;
        RECT 215.310 41.600 219.230 41.880 ;
        RECT 220.910 41.600 226.510 41.880 ;
        RECT 214.470 41.320 218.950 41.600 ;
        RECT 220.630 41.320 226.230 41.600 ;
        RECT 213.350 41.040 218.390 41.320 ;
        RECT 220.070 41.040 225.950 41.320 ;
        RECT 211.670 40.760 217.830 41.040 ;
        RECT 219.790 40.760 225.670 41.040 ;
        RECT 181.150 40.200 183.110 40.760 ;
        RECT 194.870 40.480 201.030 40.760 ;
        RECT 202.990 40.480 217.270 40.760 ;
        RECT 219.230 40.480 225.390 40.760 ;
        RECT 195.150 40.200 201.590 40.480 ;
        RECT 203.550 40.200 216.710 40.480 ;
        RECT 218.950 40.200 225.110 40.480 ;
        RECT 167.150 39.920 170.230 40.200 ;
        RECT 175.550 39.920 183.110 40.200 ;
        RECT 195.710 39.920 202.150 40.200 ;
        RECT 204.390 39.920 216.150 40.200 ;
        RECT 218.390 39.920 224.830 40.200 ;
        RECT 167.430 39.640 170.230 39.920 ;
        RECT 175.270 39.640 183.110 39.920 ;
        RECT 195.990 39.640 202.710 39.920 ;
        RECT 205.230 39.640 215.310 39.920 ;
        RECT 217.830 39.640 224.550 39.920 ;
        RECT 156.790 39.080 158.470 39.360 ;
        RECT 148.950 38.800 150.630 39.080 ;
        RECT 140.830 38.520 146.430 38.800 ;
        RECT 140.830 37.680 142.790 38.520 ;
        RECT 148.670 37.680 150.630 38.800 ;
        RECT 156.510 38.520 158.470 39.080 ;
        RECT 156.510 38.240 158.190 38.520 ;
        RECT 156.230 37.680 158.190 38.240 ;
        RECT 140.830 37.400 142.510 37.680 ;
        RECT 148.670 37.400 150.350 37.680 ;
        RECT 156.230 37.400 157.910 37.680 ;
        RECT 140.550 36.280 142.510 37.400 ;
        RECT 148.390 36.280 150.350 37.400 ;
        RECT 155.950 37.120 157.910 37.400 ;
        RECT 155.950 36.840 157.630 37.120 ;
        RECT 160.710 36.840 162.670 39.360 ;
        RECT 167.710 39.360 170.510 39.640 ;
        RECT 167.710 39.080 170.790 39.360 ;
        RECT 167.990 38.800 171.070 39.080 ;
        RECT 175.270 38.800 182.830 39.640 ;
        RECT 196.270 39.360 203.270 39.640 ;
        RECT 206.070 39.360 214.190 39.640 ;
        RECT 217.270 39.360 224.270 39.640 ;
        RECT 196.550 39.080 203.830 39.360 ;
        RECT 207.750 39.080 212.790 39.360 ;
        RECT 216.430 39.080 223.990 39.360 ;
        RECT 196.830 38.800 204.670 39.080 ;
        RECT 215.590 38.800 223.430 39.080 ;
        RECT 168.270 38.520 171.350 38.800 ;
        RECT 174.990 38.520 182.830 38.800 ;
        RECT 197.110 38.520 205.790 38.800 ;
        RECT 214.750 38.520 223.150 38.800 ;
        RECT 168.550 38.240 171.630 38.520 ;
        RECT 168.830 37.960 171.910 38.240 ;
        RECT 169.110 37.680 172.190 37.960 ;
        RECT 174.990 37.680 176.950 38.520 ;
        RECT 180.870 38.240 182.550 38.520 ;
        RECT 197.670 38.240 206.910 38.520 ;
        RECT 213.630 38.240 222.870 38.520 ;
        RECT 169.390 37.400 172.470 37.680 ;
        RECT 174.990 37.400 176.670 37.680 ;
        RECT 169.670 37.120 172.470 37.400 ;
        RECT 169.950 36.840 172.470 37.120 ;
        RECT 155.950 36.560 162.670 36.840 ;
        RECT 155.670 36.280 162.670 36.560 ;
        RECT 170.230 36.560 172.470 36.840 ;
        RECT 140.550 36.000 142.230 36.280 ;
        RECT 148.390 36.000 150.070 36.280 ;
        RECT 155.670 36.000 162.390 36.280 ;
        RECT 163.230 36.000 166.590 36.280 ;
        RECT 140.270 34.880 142.230 36.000 ;
        RECT 148.110 34.880 150.070 36.000 ;
        RECT 155.390 35.160 162.390 36.000 ;
        RECT 164.630 35.440 166.590 36.000 ;
        RECT 139.990 33.760 141.950 34.880 ;
        RECT 147.830 33.760 149.790 34.880 ;
        RECT 155.110 34.600 157.070 35.160 ;
        RECT 155.110 34.320 156.790 34.600 ;
        RECT 154.830 33.760 156.790 34.320 ;
        RECT 139.990 33.480 141.670 33.760 ;
        RECT 147.830 33.480 149.510 33.760 ;
        RECT 139.710 32.360 141.670 33.480 ;
        RECT 147.550 32.360 149.510 33.480 ;
        RECT 154.550 32.920 156.510 33.760 ;
        RECT 139.710 32.080 141.390 32.360 ;
        RECT 147.550 32.080 149.230 32.360 ;
        RECT 154.270 32.080 156.230 32.920 ;
        RECT 139.430 30.960 141.390 32.080 ;
        RECT 147.270 31.800 149.230 32.080 ;
        RECT 147.270 31.240 152.870 31.800 ;
        RECT 153.990 31.520 155.950 32.080 ;
        RECT 160.430 31.800 162.390 35.160 ;
        RECT 164.350 34.320 166.310 35.440 ;
        RECT 170.230 35.160 172.190 36.560 ;
        RECT 174.710 36.280 176.670 37.400 ;
        RECT 180.590 37.120 182.550 38.240 ;
        RECT 197.950 37.960 208.870 38.240 ;
        RECT 211.670 37.960 222.310 38.240 ;
        RECT 198.510 37.680 222.030 37.960 ;
        RECT 198.790 37.400 221.470 37.680 ;
        RECT 199.350 37.120 221.190 37.400 ;
        RECT 180.590 36.840 182.270 37.120 ;
        RECT 199.910 36.840 220.630 37.120 ;
        RECT 174.710 36.000 176.390 36.280 ;
        RECT 164.350 34.040 166.030 34.320 ;
        RECT 164.070 33.200 166.030 34.040 ;
        RECT 169.950 34.040 171.910 35.160 ;
        RECT 174.430 34.880 176.390 36.000 ;
        RECT 180.310 35.720 182.270 36.840 ;
        RECT 200.190 36.560 220.070 36.840 ;
        RECT 200.750 36.280 219.510 36.560 ;
        RECT 201.590 36.000 218.950 36.280 ;
        RECT 202.150 35.720 218.390 36.000 ;
        RECT 180.310 35.440 181.990 35.720 ;
        RECT 202.710 35.440 217.550 35.720 ;
        RECT 169.950 33.760 171.630 34.040 ;
        RECT 164.070 32.920 165.750 33.200 ;
        RECT 169.670 32.920 171.630 33.760 ;
        RECT 174.150 33.760 176.110 34.880 ;
        RECT 180.030 34.600 181.990 35.440 ;
        RECT 203.550 35.160 216.710 35.440 ;
        RECT 204.670 34.880 215.870 35.160 ;
        RECT 205.790 34.600 214.470 34.880 ;
        RECT 180.030 34.320 181.710 34.600 ;
        RECT 207.470 34.320 212.790 34.600 ;
        RECT 174.150 33.480 175.830 33.760 ;
        RECT 163.790 32.360 166.030 32.920 ;
        RECT 169.390 32.640 171.630 32.920 ;
        RECT 169.110 32.360 171.350 32.640 ;
        RECT 163.790 32.080 166.310 32.360 ;
        RECT 168.830 32.080 171.350 32.360 ;
        RECT 173.870 32.360 175.830 33.480 ;
        RECT 179.750 33.200 181.710 34.320 ;
        RECT 179.750 32.920 181.430 33.200 ;
        RECT 173.870 32.080 175.550 32.360 ;
        RECT 163.790 31.800 166.590 32.080 ;
        RECT 168.550 31.800 171.350 32.080 ;
        RECT 160.150 31.520 162.390 31.800 ;
        RECT 164.070 31.520 170.790 31.800 ;
        RECT 153.990 31.240 155.670 31.520 ;
        RECT 147.270 30.960 152.590 31.240 ;
        RECT 139.150 30.120 141.110 30.960 ;
        RECT 146.990 30.120 152.590 30.960 ;
        RECT 153.710 30.680 155.670 31.240 ;
        RECT 153.430 30.120 155.390 30.680 ;
        RECT 160.150 30.120 162.110 31.520 ;
        RECT 164.350 31.240 170.510 31.520 ;
        RECT 164.630 30.960 170.230 31.240 ;
        RECT 173.590 30.960 175.550 32.080 ;
        RECT 179.470 31.800 181.430 32.920 ;
        RECT 179.470 31.520 181.150 31.800 ;
        RECT 164.630 30.680 169.950 30.960 ;
        RECT 164.910 30.400 169.390 30.680 ;
        RECT 165.190 30.120 169.110 30.400 ;
        RECT 173.310 30.120 175.270 30.960 ;
        RECT 179.190 30.680 181.150 31.520 ;
        RECT 179.190 30.400 180.870 30.680 ;
        RECT 178.910 30.120 180.870 30.400 ;
      LAYER met3 ;
        RECT 69.070 223.300 69.830 224.480 ;
        RECT 69.470 219.220 69.830 223.300 ;
        RECT 71.830 223.270 72.590 224.450 ;
        RECT 72.290 220.700 72.590 223.270 ;
        RECT 74.620 223.260 75.380 224.440 ;
        RECT 75.070 221.090 75.380 223.260 ;
        RECT 77.380 223.220 78.140 224.400 ;
        RECT 80.120 223.220 80.880 224.400 ;
        RECT 77.840 222.000 78.140 223.220 ;
        RECT 80.570 222.650 80.880 223.220 ;
        RECT 82.900 223.170 83.980 224.350 ;
        RECT 85.650 223.170 86.410 224.350 ;
        RECT 103.870 223.340 105.040 224.010 ;
        RECT 80.570 222.320 83.360 222.650 ;
        RECT 77.840 221.700 82.730 222.000 ;
        RECT 75.070 220.790 82.100 221.090 ;
        RECT 72.280 220.310 72.590 220.700 ;
        RECT 72.280 219.920 81.480 220.310 ;
        RECT 69.470 218.860 80.880 219.220 ;
        RECT 12.460 213.330 32.200 217.740 ;
        RECT 20.960 203.250 22.160 205.440 ;
        RECT 1.000 195.080 17.070 200.820 ;
        RECT 13.030 181.860 14.560 191.150 ;
        RECT 1.000 170.760 16.520 177.210 ;
        RECT 6.000 170.750 16.520 170.760 ;
        RECT 13.270 166.240 14.550 168.580 ;
        RECT 1.000 156.970 16.530 163.410 ;
        RECT 24.420 150.080 25.230 211.770 ;
        RECT 24.420 147.750 25.730 150.080 ;
        RECT 11.930 142.070 23.490 144.800 ;
        RECT 24.420 138.550 25.230 147.750 ;
        RECT 27.070 142.030 32.200 213.330 ;
        RECT 34.160 146.650 35.760 217.740 ;
        RECT 34.160 144.870 36.190 146.650 ;
        RECT 34.170 144.850 36.190 144.870 ;
        RECT 46.760 142.030 50.360 217.740 ;
        RECT 50.990 185.170 51.780 213.660 ;
        RECT 52.970 203.450 53.610 205.830 ;
        RECT 53.000 190.440 53.640 192.820 ;
        RECT 50.990 183.140 51.810 185.170 ;
        RECT 50.990 149.090 51.780 183.140 ;
        RECT 52.980 166.420 53.620 168.800 ;
        RECT 50.990 148.410 53.060 149.090 ;
        RECT 54.510 142.030 57.880 217.740 ;
        RECT 74.470 142.030 79.600 217.740 ;
        RECT 80.570 168.980 80.880 218.860 ;
        RECT 81.180 217.740 81.480 219.920 ;
        RECT 81.800 217.740 82.100 220.790 ;
        RECT 81.180 177.330 81.490 217.740 ;
        RECT 81.800 183.730 82.110 217.740 ;
        RECT 82.420 192.260 82.730 221.700 ;
        RECT 83.050 198.290 83.360 222.320 ;
        RECT 83.670 206.520 83.980 223.170 ;
        RECT 85.830 217.740 86.260 223.170 ;
        RECT 84.300 217.440 86.260 217.740 ;
        RECT 84.300 213.000 84.610 217.440 ;
        RECT 84.300 212.030 85.420 213.000 ;
        RECT 83.670 205.650 84.650 206.520 ;
        RECT 83.050 197.680 85.020 198.290 ;
        RECT 82.410 191.240 83.520 192.260 ;
        RECT 81.800 183.070 83.190 183.730 ;
        RECT 81.180 176.980 84.800 177.330 ;
        RECT 80.570 168.620 84.740 168.980 ;
        RECT 83.780 168.100 84.740 168.620 ;
        RECT 86.480 142.040 89.080 216.710 ;
        RECT 93.850 214.430 94.240 215.410 ;
        RECT 93.850 213.940 95.100 214.430 ;
        RECT 90.260 194.090 90.610 212.580 ;
        RECT 92.270 203.960 92.650 203.970 ;
        RECT 93.820 203.960 94.250 204.920 ;
        RECT 92.270 203.540 94.250 203.960 ;
        RECT 90.050 193.460 90.850 194.090 ;
        RECT 92.270 175.260 92.650 203.540 ;
        RECT 94.710 202.830 95.100 213.940 ;
        RECT 96.680 207.500 97.060 213.900 ;
        RECT 97.870 206.970 98.310 212.730 ;
        RECT 93.070 202.510 95.100 202.830 ;
        RECT 93.070 185.260 93.460 202.510 ;
        RECT 91.360 174.840 92.650 175.260 ;
        RECT 93.850 170.480 94.220 199.880 ;
        RECT 92.720 170.040 94.220 170.480 ;
        RECT 95.550 142.040 98.500 202.530 ;
        RECT 99.140 200.340 99.510 208.240 ;
        RECT 100.470 142.040 103.210 216.710 ;
        RECT 104.680 213.490 105.040 223.340 ;
        RECT 105.680 222.240 107.270 222.930 ;
        RECT 104.630 212.320 105.100 213.490 ;
        RECT 105.680 207.320 106.000 222.240 ;
        RECT 107.150 221.060 108.590 221.480 ;
        RECT 105.610 206.150 106.080 207.320 ;
        RECT 107.150 198.930 107.510 221.060 ;
        RECT 107.100 197.760 107.570 198.930 ;
        RECT 23.900 132.410 25.960 138.550 ;
      LAYER met4 ;
        RECT 69.310 224.480 69.610 224.760 ;
        RECT 69.070 223.300 69.830 224.480 ;
        RECT 72.070 224.450 72.370 224.760 ;
        RECT 71.830 223.270 72.590 224.450 ;
        RECT 74.830 224.440 75.130 224.760 ;
        RECT 74.620 223.260 75.380 224.440 ;
        RECT 77.590 224.400 77.890 224.760 ;
        RECT 80.350 224.400 80.650 224.760 ;
        RECT 77.380 223.220 78.140 224.400 ;
        RECT 80.120 223.220 80.880 224.400 ;
        RECT 83.110 224.350 83.410 224.760 ;
        RECT 85.870 224.350 86.170 224.760 ;
        RECT 82.900 223.170 83.660 224.350 ;
        RECT 85.650 223.170 86.410 224.350 ;
        RECT 88.630 221.480 88.930 224.760 ;
        RECT 91.390 222.580 91.690 224.760 ;
        RECT 94.150 223.710 94.450 224.760 ;
        RECT 103.870 223.710 105.040 224.010 ;
        RECT 94.150 223.340 105.040 223.710 ;
        RECT 105.680 222.580 107.270 222.930 ;
        RECT 91.390 222.240 107.270 222.580 ;
        RECT 88.630 221.060 108.590 221.480 ;
        RECT 6.000 213.330 103.210 217.740 ;
        RECT 20.960 205.050 22.160 205.440 ;
        RECT 52.970 205.050 53.610 205.830 ;
        RECT 20.960 204.300 53.610 205.050 ;
        RECT 20.960 203.250 22.160 204.300 ;
        RECT 52.970 203.450 53.610 204.300 ;
        RECT 8.390 195.080 102.980 200.820 ;
        RECT 53.000 191.150 53.640 192.820 ;
        RECT 13.030 190.440 53.640 191.150 ;
        RECT 13.030 189.780 14.560 190.440 ;
        RECT 6.000 180.550 103.210 185.990 ;
        RECT 8.470 170.750 103.100 177.230 ;
        RECT 13.270 168.050 14.560 168.600 ;
        RECT 52.980 168.050 53.620 168.800 ;
        RECT 13.270 167.200 53.620 168.050 ;
        RECT 13.270 166.250 14.560 167.200 ;
        RECT 52.980 166.420 53.620 167.200 ;
        RECT 8.400 156.980 103.200 163.420 ;
        RECT 6.000 148.770 103.220 153.780 ;
        RECT 11.930 142.070 23.490 144.800 ;
        RECT 16.630 6.500 18.050 142.070 ;
        RECT 23.900 132.410 25.960 138.550 ;
        RECT 24.410 11.050 25.460 132.410 ;
        RECT 24.340 9.850 152.710 11.050 ;
        RECT 16.630 5.300 133.390 6.500 ;
        RECT 16.630 5.290 18.440 5.300 ;
        RECT 132.490 1.000 133.390 5.300 ;
        RECT 151.810 1.000 152.710 9.850 ;
  END
END tt_um_tinyflash
END LIBRARY

