magic
tech sky130A
magscale 1 2
timestamp 1762640459
<< pwell >>
rect -739 -1155 739 1155
<< psubdiff >>
rect -703 1085 -607 1119
rect 607 1085 703 1119
rect -703 -1085 -669 1085
rect 669 -1085 703 1085
rect -703 -1119 -607 -1085
rect 607 -1119 703 -1085
<< psubdiffcont >>
rect -607 1085 607 1119
rect -607 -1119 607 -1085
<< xpolycontact >>
rect -573 557 573 989
rect -573 -989 573 -557
<< xpolyres >>
rect -573 -557 573 557
<< locali >>
rect -703 1085 -607 1119
rect 607 1085 703 1119
rect -703 -1085 -669 1085
rect 669 -1085 703 1085
rect -703 -1119 -607 -1085
rect 607 -1119 703 -1085
<< viali >>
rect -557 574 557 971
rect -557 -971 557 -574
<< metal1 >>
rect -569 971 569 977
rect -569 574 -557 971
rect 557 574 569 971
rect -569 568 569 574
rect -569 -574 569 -568
rect -569 -971 -557 -574
rect 557 -971 569 -574
rect -569 -977 569 -971
<< labels >>
rlabel psubdiffcont 0 -1102 0 -1102 0 B
port 28 nsew
rlabel xpolycontact 0 954 0 954 0 R1
port 29 nsew
rlabel xpolycontact 0 -954 0 -954 0 R2
port 30 nsew
<< properties >>
string FIXED_BBOX -686 -1102 686 1102
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 5.73 m 1 nx 1 wmin 5.730 lmin 0.50 class resistor rho 2000 val 2.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 doports 1 mult 1
<< end >>
