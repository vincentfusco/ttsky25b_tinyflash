magic
tech sky130A
timestamp 1762644791
<< pwell >>
rect -153 -641 153 641
<< psubdiff >>
rect -135 606 -87 623
rect 87 606 135 623
rect -135 -606 -118 606
rect 118 -606 135 606
rect -135 -623 -87 -606
rect 87 -623 135 -606
<< psubdiffcont >>
rect -87 606 87 623
rect -87 -623 87 -606
<< xpolycontact >>
rect -70 342 70 558
rect -70 -558 70 -342
<< xpolyres >>
rect -70 -342 70 342
<< locali >>
rect -135 606 -87 623
rect 87 606 135 623
rect -135 -606 -118 606
rect 118 -606 135 606
rect -135 -623 -87 -606
rect 87 -623 135 -606
<< viali >>
rect -62 350 62 549
rect -62 -549 62 -350
<< metal1 >>
rect -65 549 65 555
rect -65 350 -62 549
rect 62 350 65 549
rect -65 344 65 350
rect -65 -350 65 -344
rect -65 -549 -62 -350
rect 62 -549 65 -350
rect -65 -555 65 -549
<< labels >>
rlabel psubdiffcont 0 -614 0 -614 0 B
port 10 nsew
rlabel xpolycontact 0 540 0 540 0 R1
port 11 nsew
rlabel xpolycontact 0 -540 0 -540 0 R2
port 12 nsew
<< properties >>
string FIXED_BBOX -127 -614 127 614
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 7.0 m 1 nx 1 wmin 1.410 lmin 0.50 class resistor rho 2000 val 10.196k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 doports 1 mult 1
<< end >>
