* NGSPICE file created from res_ladder_vref_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_5p73_JT48NU B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_5p73 l=5.73
C0 R2 R1 0.06813f
C1 R2 B 1.74197f
C2 R1 B 1.74197f
.ends

.subckt res_ladder_vref_extracted ref0 ref1 ref2 ref3 ref4 ref5 ref6 vref vss
XXR1 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR2 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR10 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR3 vss ref6 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR4 vss ref4 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR5 vss ref4 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR6 vss ref2 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR7 vss ref2 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR8 vss ref0 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR9 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
R0 ref6.n0 ref6 2.13017
R1 ref6.n1 ref6 2.13017
R2 ref6.n2 ref6 2.13017
R3 ref6.n2 ref6.n1 0.397491
R4 ref6.n1 ref6.n0 0.397491
R5 ref6 ref6.n2 0.166299
R6 ref6.n0 ref6 0.166299
R7 vref.n0 vref 2.51601
R8 vref.n0 vref 2.11902
R9 vref vref.n1 1.37411
R10 vref.n1 vref 0.831056
R11 vref.n1 vref 0.774111
R12 vref.n1 vref 0.231056
R13 vref vref.n0 0.188289
R14 vref.n1 vref 0.0135208
R15 vref.n1 vref 0.0135208
R16 vss.n108 vss.n3 10261.4
R17 vss.n40 vss.n39 10261.4
R18 vss.n101 vss.n5 6385.12
R19 vss.n101 vss.n2 6385.12
R20 vss.n94 vss.n7 6385.12
R21 vss.n94 vss.n9 6385.12
R22 vss.n87 vss.n13 6385.12
R23 vss.n87 vss.n11 6385.12
R24 vss.n80 vss.n15 6385.12
R25 vss.n80 vss.n17 6385.12
R26 vss.n73 vss.n21 6385.12
R27 vss.n73 vss.n19 6385.12
R28 vss.n66 vss.n23 6385.12
R29 vss.n66 vss.n25 6385.12
R30 vss.n59 vss.n29 6385.12
R31 vss.n59 vss.n27 6385.12
R32 vss.n52 vss.n31 6385.12
R33 vss.n52 vss.n33 6385.12
R34 vss.n45 vss.n37 6385.12
R35 vss.n45 vss.n35 6385.12
R36 vss.n108 vss.n2 3876.26
R37 vss.n99 vss.n7 3876.26
R38 vss.n99 vss.n5 3876.26
R39 vss.n105 vss.n5 3876.26
R40 vss.n93 vss.n11 3876.26
R41 vss.n93 vss.n9 3876.26
R42 vss.n97 vss.n9 3876.26
R43 vss.n97 vss.n2 3876.26
R44 vss.n85 vss.n15 3876.26
R45 vss.n85 vss.n13 3876.26
R46 vss.n91 vss.n13 3876.26
R47 vss.n91 vss.n7 3876.26
R48 vss.n79 vss.n19 3876.26
R49 vss.n79 vss.n17 3876.26
R50 vss.n83 vss.n17 3876.26
R51 vss.n83 vss.n11 3876.26
R52 vss.n71 vss.n23 3876.26
R53 vss.n71 vss.n21 3876.26
R54 vss.n77 vss.n21 3876.26
R55 vss.n77 vss.n15 3876.26
R56 vss.n65 vss.n27 3876.26
R57 vss.n65 vss.n25 3876.26
R58 vss.n69 vss.n25 3876.26
R59 vss.n69 vss.n19 3876.26
R60 vss.n57 vss.n31 3876.26
R61 vss.n57 vss.n29 3876.26
R62 vss.n63 vss.n29 3876.26
R63 vss.n63 vss.n23 3876.26
R64 vss.n51 vss.n35 3876.26
R65 vss.n51 vss.n33 3876.26
R66 vss.n55 vss.n33 3876.26
R67 vss.n55 vss.n27 3876.26
R68 vss.n43 vss.n37 3876.26
R69 vss.n49 vss.n37 3876.26
R70 vss.n49 vss.n31 3876.26
R71 vss.n40 vss.n35 3876.26
R72 vss.n41 vss.n36 1306.67
R73 vss.n50 vss.n36 1306.67
R74 vss.n50 vss.n32 1306.67
R75 vss.n56 vss.n32 1306.67
R76 vss.n56 vss.n28 1306.67
R77 vss.n64 vss.n28 1306.67
R78 vss.n64 vss.n24 1306.67
R79 vss.n70 vss.n24 1306.67
R80 vss.n70 vss.n20 1306.67
R81 vss.n78 vss.n20 1306.67
R82 vss.n78 vss.n16 1306.67
R83 vss.n84 vss.n16 1306.67
R84 vss.n84 vss.n12 1306.67
R85 vss.n92 vss.n12 1306.67
R86 vss.n92 vss.n8 1306.67
R87 vss.n98 vss.n8 1306.67
R88 vss.n98 vss.n4 1306.67
R89 vss.n107 vss.n4 1306.67
R90 vss.n106 vss.n3 1171.11
R91 vss.n42 vss.n39 1171.11
R92 vss vss.n38 666.73
R93 vss.n44 vss.n38 666.73
R94 vss.n104 vss.n0 621.553
R95 vss.n109 vss 619.196
R96 vss.n47 vss.n46 414.872
R97 vss.n46 vss.n34 414.872
R98 vss.n53 vss.n30 414.872
R99 vss.n54 vss.n53 414.872
R100 vss.n61 vss.n60 414.872
R101 vss.n60 vss.n26 414.872
R102 vss.n67 vss.n22 414.872
R103 vss.n68 vss.n67 414.872
R104 vss.n75 vss.n74 414.872
R105 vss.n74 vss.n18 414.872
R106 vss.n81 vss.n14 414.872
R107 vss.n82 vss.n81 414.872
R108 vss.n89 vss.n88 414.872
R109 vss.n88 vss.n10 414.872
R110 vss.n95 vss.n6 414.872
R111 vss.n96 vss.n95 414.872
R112 vss.n103 vss.n102 414.872
R113 vss.n102 vss.n1 414.872
R114 vss vss.n34 251.859
R115 vss.n47 vss.n44 251.859
R116 vss.n48 vss.n47 251.859
R117 vss.n48 vss.n30 251.859
R118 vss vss.n34 251.859
R119 vss.n54 vss 251.859
R120 vss vss.n54 251.859
R121 vss vss.n26 251.859
R122 vss.n58 vss.n30 251.859
R123 vss.n61 vss.n58 251.859
R124 vss.n62 vss.n61 251.859
R125 vss.n62 vss.n22 251.859
R126 vss vss.n26 251.859
R127 vss.n68 vss 251.859
R128 vss vss.n68 251.859
R129 vss vss.n18 251.859
R130 vss.n72 vss.n22 251.859
R131 vss.n75 vss.n72 251.859
R132 vss.n76 vss.n75 251.859
R133 vss.n76 vss.n14 251.859
R134 vss vss.n18 251.859
R135 vss.n82 vss 251.859
R136 vss vss.n82 251.859
R137 vss vss.n10 251.859
R138 vss.n86 vss.n14 251.859
R139 vss.n89 vss.n86 251.859
R140 vss.n90 vss.n89 251.859
R141 vss.n90 vss.n6 251.859
R142 vss vss.n10 251.859
R143 vss.n96 vss 251.859
R144 vss vss.n96 251.859
R145 vss vss.n1 251.859
R146 vss.n100 vss.n6 251.859
R147 vss.n103 vss.n100 251.859
R148 vss.n104 vss.n103 251.859
R149 vss vss.n1 251.859
R150 vss.n40 vss 32.5005
R151 vss.n41 vss.n40 32.5005
R152 vss.n44 vss.n43 32.5005
R153 vss.n49 vss.n48 32.5005
R154 vss.n50 vss.n49 32.5005
R155 vss vss.n51 32.5005
R156 vss.n51 vss.n50 32.5005
R157 vss.n55 vss 32.5005
R158 vss.n56 vss.n55 32.5005
R159 vss.n58 vss.n57 32.5005
R160 vss.n57 vss.n56 32.5005
R161 vss.n63 vss.n62 32.5005
R162 vss.n64 vss.n63 32.5005
R163 vss vss.n65 32.5005
R164 vss.n65 vss.n64 32.5005
R165 vss.n69 vss 32.5005
R166 vss.n70 vss.n69 32.5005
R167 vss.n72 vss.n71 32.5005
R168 vss.n71 vss.n70 32.5005
R169 vss.n77 vss.n76 32.5005
R170 vss.n78 vss.n77 32.5005
R171 vss vss.n79 32.5005
R172 vss.n79 vss.n78 32.5005
R173 vss.n83 vss 32.5005
R174 vss.n84 vss.n83 32.5005
R175 vss.n86 vss.n85 32.5005
R176 vss.n85 vss.n84 32.5005
R177 vss.n91 vss.n90 32.5005
R178 vss.n92 vss.n91 32.5005
R179 vss vss.n93 32.5005
R180 vss.n93 vss.n92 32.5005
R181 vss.n97 vss 32.5005
R182 vss.n98 vss.n97 32.5005
R183 vss.n100 vss.n99 32.5005
R184 vss.n99 vss.n98 32.5005
R185 vss.n105 vss.n104 32.5005
R186 vss vss.n108 32.5005
R187 vss.n108 vss.n107 32.5005
R188 vss.n106 vss.n105 28.701
R189 vss.n43 vss.n42 28.701
R190 vss.n39 vss.n38 19.5005
R191 vss.n46 vss.n45 19.5005
R192 vss.n45 vss.n36 19.5005
R193 vss.n53 vss.n52 19.5005
R194 vss.n52 vss.n32 19.5005
R195 vss.n60 vss.n59 19.5005
R196 vss.n59 vss.n28 19.5005
R197 vss.n67 vss.n66 19.5005
R198 vss.n66 vss.n24 19.5005
R199 vss.n74 vss.n73 19.5005
R200 vss.n73 vss.n20 19.5005
R201 vss.n81 vss.n80 19.5005
R202 vss.n80 vss.n16 19.5005
R203 vss.n88 vss.n87 19.5005
R204 vss.n87 vss.n12 19.5005
R205 vss.n95 vss.n94 19.5005
R206 vss.n94 vss.n8 19.5005
R207 vss.n102 vss.n101 19.5005
R208 vss.n101 vss.n4 19.5005
R209 vss.n3 vss.n0 19.5005
R210 vss.n42 vss.n41 3.71014
R211 vss.n107 vss.n106 3.71014
R212 vss.n111 vss 2.51601
R213 vss.n109 vss.n0 2.35839
R214 vss.n111 vss 2.11902
R215 vss vss.n112 1.37411
R216 vss.n112 vss 0.831056
R217 vss.n112 vss.n110 0.764389
R218 vss.n110 vss.n109 0.3005
R219 vss.n112 vss 0.231056
R220 vss.n112 vss.n111 0.20131
R221 vss.n110 vss 0.0102222
R222 vss.n112 vss 0.00426157
R223 ref0.n0 ref0 2.13017
R224 ref0.n1 ref0 2.13017
R225 ref0.n2 ref0 2.13017
R226 ref0.n2 ref0.n1 0.397491
R227 ref0.n1 ref0.n0 0.397491
R228 ref0 ref0.n2 0.166299
R229 ref0.n0 ref0 0.166299
R230 ref5.n1 ref5 2.11902
R231 ref5.n0 ref5 2.11902
R232 ref5.n1 ref5.n0 0.397491
R233 ref5 ref5.n1 0.166299
R234 ref5.n0 ref5 0.166299
R235 ref4.n0 ref4 2.13017
R236 ref4.n1 ref4 2.13017
R237 ref4.n1 ref4.n0 0.397491
R238 ref4 ref4.n1 0.166299
R239 ref4.n0 ref4 0.166299
R240 ref3.n1 ref3 2.11902
R241 ref3.n0 ref3 2.11902
R242 ref3.n1 ref3.n0 0.397491
R243 ref3 ref3.n1 0.166299
R244 ref3.n0 ref3 0.166299
R245 ref2.n0 ref2 2.13017
R246 ref2.n1 ref2 2.13017
R247 ref2.n1 ref2.n0 0.397491
R248 ref2 ref2.n1 0.166299
R249 ref2.n0 ref2 0.166299
R250 ref1.n1 ref1 2.11902
R251 ref1.n0 ref1 2.11902
R252 ref1.n1 ref1.n0 0.397491
R253 ref1 ref1.n1 0.166299
R254 ref1.n0 ref1 0.166299
C0 ref2 ref3 0
C1 ref6 ref5 0
C2 ref5 ref4 0
C3 vref ref6 0.16095f
C4 ref2 ref1 0
C5 ref5 ref3 0.06887f
C6 ref2 ref0 0.06887f
C7 ref3 ref1 0.06887f
C8 vref ref5 0.06887f
C9 ref6 ref4 0.06887f
C10 ref2 ref4 0.06887f
C11 ref1 ref0 0
C12 ref4 ref3 0
C13 ref0 vss 5.32418f
C14 ref1 vss 3.4889f
C15 ref2 vss 3.42003f
C16 ref3 vss 3.42003f
C17 ref4 vss 3.42003f
C18 ref5 vss 3.42003f
C19 ref6 vss 5.161f
C20 vref vss 4.57377f
.ends

