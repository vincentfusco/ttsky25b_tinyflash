VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO flashADC_3bit
  CLASS BLOCK ;
  FOREIGN flashADC_3bit ;
  ORIGIN 15.350 57.070 ;
  SIZE 93.120 BY 80.030 ;
  PIN vin
    ANTENNAGATEAREA 97.950996 ;
    PORT
      LAYER met3 ;
        RECT -2.870 -56.220 -2.060 -44.100 ;
    END
  END vin
  PIN vref
    PORT
      LAYER met1 ;
        RECT -15.350 -53.890 -3.800 -53.440 ;
    END
  END vref
  PIN dout0
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met1 ;
        RECT 76.340 14.080 76.800 14.480 ;
    END
  END dout0
  PIN dout1
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met1 ;
        RECT 76.340 7.880 76.800 8.280 ;
    END
  END dout1
  PIN dout2
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met1 ;
        RECT 76.340 -0.500 76.800 -0.100 ;
    END
  END dout2
  PIN d0
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met3 ;
        RECT 57.010 14.590 57.320 19.500 ;
    END
  END d0
  PIN d1
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met3 ;
        RECT 56.380 8.140 56.690 19.500 ;
    END
  END d1
  PIN d2
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met3 ;
        RECT 55.760 -0.560 56.070 19.500 ;
    END
  END d2
  PIN d3
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met3 ;
        RECT 55.130 -6.620 55.440 19.500 ;
    END
  END d3
  PIN d4
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met3 ;
        RECT 54.510 -14.550 54.820 19.500 ;
    END
  END d4
  PIN d5
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met3 ;
        RECT 53.890 -21.260 54.200 -20.920 ;
    END
  END d5
  PIN d6
    ANTENNAGATEAREA 0.450000 ;
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER met3 ;
        RECT 53.280 -29.620 53.590 19.500 ;
    END
  END d6
  PIN vdd
    ANTENNADIFFAREA 283.898590 ;
    PORT
      LAYER met3 ;
        RECT 27.220 19.130 30.590 19.500 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 265.982391 ;
    PORT
      LAYER met3 ;
        RECT -0.220 0.940 4.910 19.500 ;
    END
  END vss
  OBS
      LAYER pwell ;
        RECT -15.350 18.470 77.770 22.960 ;
        RECT -15.350 5.350 -0.220 18.470 ;
      LAYER nwell ;
        RECT -0.220 5.350 77.770 18.470 ;
      LAYER pwell ;
        RECT -15.350 -0.300 57.890 5.350 ;
      LAYER nwell ;
        RECT 57.890 -0.300 77.770 5.350 ;
      LAYER pwell ;
        RECT -15.350 -3.400 77.770 -0.300 ;
        RECT -15.350 -3.690 73.380 -3.400 ;
      LAYER nwell ;
        RECT 73.380 -3.690 77.770 -3.400 ;
      LAYER pwell ;
        RECT -15.350 -5.430 77.770 -3.690 ;
        RECT -15.350 -31.670 -0.220 -5.430 ;
      LAYER nwell ;
        RECT -0.220 -31.670 77.770 -5.430 ;
      LAYER pwell ;
        RECT -15.350 -42.450 77.770 -31.670 ;
        RECT -15.350 -52.770 23.520 -42.450 ;
      LAYER nwell ;
        RECT 23.520 -52.770 77.770 -42.450 ;
      LAYER pwell ;
        RECT -15.350 -55.570 10.690 -52.770 ;
      LAYER nwell ;
        RECT 10.690 -55.570 77.770 -52.770 ;
      LAYER pwell ;
        RECT -15.350 -57.070 77.770 -55.570 ;
      LAYER li1 ;
        RECT -15.170 -55.390 76.670 18.330 ;
      LAYER met1 ;
        RECT -15.350 14.760 76.850 19.500 ;
        RECT -15.350 13.800 76.060 14.760 ;
        RECT -15.350 8.560 76.850 13.800 ;
        RECT -15.350 7.600 76.060 8.560 ;
        RECT -15.350 0.180 76.850 7.600 ;
        RECT -15.350 -0.780 76.060 0.180 ;
        RECT -15.350 -53.160 76.850 -0.780 ;
        RECT -15.350 -54.170 -3.800 -53.890 ;
        RECT -3.520 -54.170 76.850 -53.160 ;
        RECT -15.350 -56.210 76.850 -54.170 ;
      LAYER met2 ;
        RECT -14.830 -56.020 76.850 19.280 ;
      LAYER met3 ;
        RECT -14.830 0.540 -0.620 19.500 ;
        RECT 5.310 18.730 26.820 19.500 ;
        RECT 30.990 18.730 52.880 19.500 ;
        RECT 5.310 0.540 52.880 18.730 ;
        RECT -14.830 -30.020 52.880 0.540 ;
        RECT 53.990 -14.950 54.110 19.500 ;
        RECT 57.720 14.190 75.920 19.500 ;
        RECT 57.090 7.740 75.920 14.190 ;
        RECT 56.470 -0.960 75.920 7.740 ;
        RECT 55.840 -7.020 75.920 -0.960 ;
        RECT 55.220 -14.950 75.920 -7.020 ;
        RECT 53.990 -20.520 75.920 -14.950 ;
        RECT 54.600 -21.660 75.920 -20.520 ;
        RECT 53.990 -30.020 75.920 -21.660 ;
        RECT -14.830 -43.700 75.920 -30.020 ;
        RECT -14.830 -56.210 -3.270 -43.700 ;
        RECT -1.660 -56.210 75.920 -43.700 ;
      LAYER met4 ;
        RECT -14.260 -31.990 26.350 7.590 ;
  END
END flashADC_3bit
END LIBRARY

