magic
tech sky130A
timestamp 1762640459
<< pwell >>
rect 10561 20615 10604 20732
rect 10710 19776 10753 19893
<< metal1 >>
rect 10463 21342 10510 21349
rect 10463 21272 10471 21342
rect 10401 21238 10471 21272
rect 10503 21238 10510 21342
rect 10401 21232 10510 21238
rect 10561 20725 10608 20732
rect 10561 20652 10569 20725
rect 10363 20621 10569 20652
rect 10601 20621 10608 20725
rect 10363 20612 10608 20621
rect 10710 19886 10757 19893
rect 10710 19814 10718 19886
rect 10363 19782 10718 19814
rect 10750 19782 10757 19886
rect 10363 19774 10757 19782
rect 1193 14429 2349 14480
rect 1193 14250 1222 14429
rect 2301 14250 2349 14429
rect 1193 14207 2349 14250
<< via1 >>
rect 10471 21238 10503 21342
rect 10569 20621 10601 20725
rect 10718 19782 10750 19886
rect 1222 14250 2301 14429
<< metal2 >>
rect 10463 21342 10510 21349
rect 10463 21238 10471 21342
rect 10503 21238 10510 21342
rect 10463 21232 10510 21238
rect 10561 20725 10608 20732
rect 10561 20621 10569 20725
rect 10601 20621 10608 20725
rect 10561 20615 10608 20621
rect 10710 19886 10757 19893
rect 10710 19782 10718 19886
rect 10750 19782 10757 19886
rect 10710 19776 10757 19782
rect 1193 14429 2349 14480
rect 1193 14250 1222 14429
rect 2301 14250 2349 14429
rect 1193 14207 2349 14250
<< via2 >>
rect 10471 21238 10503 21342
rect 10569 20621 10601 20725
rect 10718 19782 10750 19886
rect 1222 14250 2301 14429
<< metal3 >>
rect 6907 22438 6983 22448
rect 6907 22343 6922 22438
rect 6968 22343 6983 22438
rect 6907 22330 6983 22343
rect 6947 21922 6983 22330
rect 7183 22435 7259 22445
rect 7183 22340 7198 22435
rect 7244 22340 7259 22435
rect 7183 22327 7259 22340
rect 7229 22070 7259 22327
rect 7462 22434 7538 22444
rect 7462 22339 7477 22434
rect 7523 22339 7538 22434
rect 7462 22326 7538 22339
rect 7507 22109 7538 22326
rect 7738 22430 7814 22440
rect 7738 22335 7753 22430
rect 7799 22335 7814 22430
rect 7738 22322 7814 22335
rect 8012 22430 8088 22440
rect 8012 22335 8027 22430
rect 8073 22335 8088 22430
rect 8012 22322 8088 22335
rect 7784 22200 7814 22322
rect 8057 22265 8088 22322
rect 8290 22425 8398 22435
rect 8290 22330 8305 22425
rect 8351 22330 8398 22425
rect 8290 22317 8398 22330
rect 8565 22425 8641 22435
rect 8565 22330 8580 22425
rect 8626 22330 8641 22425
rect 10387 22388 10504 22401
rect 10387 22350 10401 22388
rect 10490 22350 10504 22388
rect 10387 22334 10504 22350
rect 8565 22317 8641 22330
rect 8057 22232 8336 22265
rect 7784 22170 8273 22200
rect 7507 22079 8210 22109
rect 7228 22031 7259 22070
rect 7228 21992 8148 22031
rect 6947 21886 8088 21922
rect 8057 21738 8088 21886
rect 8118 21722 8148 21992
rect 8180 21761 8210 22079
rect 8242 21754 8273 22170
rect 8305 21728 8336 22232
rect 8367 21737 8398 22317
rect 8583 21774 8626 22317
rect 8430 21744 8626 21774
rect 10468 21349 10504 22334
rect 10568 22278 10727 22293
rect 10568 22237 10577 22278
rect 10712 22237 10727 22278
rect 10568 22224 10727 22237
rect 10463 21342 10510 21349
rect 10463 21238 10471 21342
rect 10503 21238 10510 21342
rect 10463 21232 10510 21238
rect 10568 20732 10600 22224
rect 10715 22144 10859 22148
rect 10715 22112 10720 22144
rect 10850 22112 10859 22144
rect 10715 22106 10859 22112
rect 10561 20725 10608 20732
rect 10561 20621 10569 20725
rect 10601 20621 10608 20725
rect 10561 20615 10608 20621
rect 100 20025 1707 20082
rect 100 19565 142 20025
rect 243 19994 1707 20025
rect 243 19596 1008 19994
rect 1647 19596 1707 19994
rect 243 19565 1707 19596
rect 100 19508 1707 19565
rect 10715 19893 10751 22106
rect 10710 19886 10757 19893
rect 10710 19782 10718 19886
rect 10750 19782 10757 19886
rect 10710 19776 10757 19782
rect 100 17661 1652 17721
rect 100 17112 143 17661
rect 255 17587 1652 17661
rect 255 17207 950 17587
rect 1526 17207 1652 17587
rect 255 17112 1652 17207
rect 100 17076 1652 17112
rect 600 17075 1652 17076
rect 100 16270 1653 16341
rect 100 15774 130 16270
rect 270 15774 882 16270
rect 1523 15774 1653 16270
rect 100 15697 1653 15774
rect 1193 14429 2349 14480
rect 1193 14250 1222 14429
rect 2301 14250 2349 14429
rect 1193 14207 2349 14250
rect 2442 13855 2523 14240
rect 2390 13811 2596 13855
rect 2390 13290 2422 13811
rect 2562 13290 2596 13811
rect 2390 13241 2596 13290
<< via3 >>
rect 6922 22343 6968 22438
rect 7198 22340 7244 22435
rect 7477 22339 7523 22434
rect 7753 22335 7799 22430
rect 8027 22335 8073 22430
rect 8305 22330 8351 22425
rect 8580 22330 8626 22425
rect 10401 22350 10490 22388
rect 1327 21420 3091 21681
rect 4713 21366 5001 21741
rect 10084 21369 10273 21631
rect 10577 22237 10712 22278
rect 10720 22112 10850 22144
rect 142 19565 243 20025
rect 1008 19596 1647 19994
rect 5502 19561 5727 20010
rect 7528 19581 7869 20000
rect 8699 19552 8847 20054
rect 9627 19547 9775 20049
rect 2791 18138 3133 18508
rect 4743 18131 4965 18523
rect 10119 18126 10265 18507
rect 143 17112 255 17661
rect 950 17207 1526 17587
rect 5503 17137 5708 17632
rect 7513 17141 7859 17622
rect 8694 17132 8842 17634
rect 9637 17134 9785 17636
rect 130 15774 270 16270
rect 882 15774 1523 16270
rect 5515 15756 5705 16249
rect 7542 15796 7860 16232
rect 8701 15763 8849 16265
rect 9629 15763 9777 16265
rect 2797 14945 3133 15295
rect 4753 14950 4945 15302
rect 10113 14946 10259 15327
rect 1222 14250 2301 14429
rect 2422 13290 2562 13811
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22448 6961 22576
rect 6907 22438 6983 22448
rect 7207 22445 7237 22576
rect 6907 22343 6922 22438
rect 6968 22343 6983 22438
rect 6907 22330 6983 22343
rect 7183 22435 7259 22445
rect 7483 22444 7513 22576
rect 7183 22340 7198 22435
rect 7244 22340 7259 22435
rect 7183 22327 7259 22340
rect 7462 22434 7538 22444
rect 7759 22440 7789 22576
rect 8035 22440 8065 22576
rect 7462 22339 7477 22434
rect 7523 22339 7538 22434
rect 7462 22326 7538 22339
rect 7738 22430 7814 22440
rect 7738 22335 7753 22430
rect 7799 22335 7814 22430
rect 7738 22322 7814 22335
rect 8012 22430 8088 22440
rect 8311 22435 8341 22576
rect 8587 22435 8617 22576
rect 8012 22335 8027 22430
rect 8073 22335 8088 22430
rect 8012 22322 8088 22335
rect 8290 22425 8366 22435
rect 8290 22330 8305 22425
rect 8351 22330 8366 22425
rect 8290 22317 8366 22330
rect 8565 22425 8641 22435
rect 8565 22330 8580 22425
rect 8626 22330 8641 22425
rect 8565 22317 8641 22330
rect 8863 22148 8893 22576
rect 9139 22258 9169 22576
rect 9415 22371 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 10387 22388 10504 22401
rect 10387 22371 10401 22388
rect 9415 22350 10401 22371
rect 10490 22350 10504 22388
rect 9415 22334 10504 22350
rect 10568 22278 10727 22293
rect 10568 22258 10577 22278
rect 9139 22237 10577 22258
rect 10712 22237 10727 22278
rect 9139 22224 10727 22237
rect 8863 22144 10859 22148
rect 8863 22112 10720 22144
rect 10850 22112 10859 22144
rect 8863 22106 10859 22112
rect 100 20025 300 22076
rect 100 19565 142 20025
rect 243 19565 300 20025
rect 100 17661 300 19565
rect 100 17112 143 17661
rect 255 17112 300 17661
rect 100 16270 300 17112
rect 100 15774 130 16270
rect 270 15774 300 16270
rect 100 500 300 15774
rect 400 21774 600 22076
rect 400 21741 10321 21774
rect 400 21681 4713 21741
rect 400 21420 1327 21681
rect 3091 21420 4713 21681
rect 400 21366 4713 21420
rect 5001 21631 10321 21741
rect 5001 21369 10084 21631
rect 10273 21369 10321 21631
rect 5001 21366 10321 21369
rect 400 21333 10321 21366
rect 400 18599 600 21333
rect 839 20054 10298 20082
rect 839 20010 8699 20054
rect 839 19994 5502 20010
rect 839 19596 1008 19994
rect 1647 19596 5502 19994
rect 839 19561 5502 19596
rect 5727 20000 8699 20010
rect 5727 19581 7528 20000
rect 7869 19581 8699 20000
rect 5727 19561 8699 19581
rect 839 19552 8699 19561
rect 8847 20049 10298 20054
rect 8847 19552 9627 20049
rect 839 19547 9627 19552
rect 9775 19547 10298 20049
rect 839 19508 10298 19547
rect 400 18523 10321 18599
rect 400 18508 4743 18523
rect 400 18138 2791 18508
rect 3133 18138 4743 18508
rect 400 18131 4743 18138
rect 4965 18507 10321 18523
rect 4965 18131 10119 18507
rect 400 18126 10119 18131
rect 10265 18126 10321 18507
rect 400 18055 10321 18126
rect 400 15378 600 18055
rect 847 17636 10310 17723
rect 847 17634 9637 17636
rect 847 17632 8694 17634
rect 847 17587 5503 17632
rect 847 17207 950 17587
rect 1526 17207 5503 17587
rect 847 17137 5503 17207
rect 5708 17622 8694 17632
rect 5708 17141 7513 17622
rect 7859 17141 8694 17622
rect 5708 17137 8694 17141
rect 847 17132 8694 17137
rect 8842 17134 9637 17634
rect 9785 17134 10310 17636
rect 8842 17132 10310 17134
rect 847 17075 10310 17132
rect 840 16270 10320 16342
rect 840 15774 882 16270
rect 1523 16265 10320 16270
rect 1523 16249 8701 16265
rect 1523 15774 5515 16249
rect 840 15756 5515 15774
rect 5705 16232 8701 16249
rect 5705 15796 7542 16232
rect 7860 15796 8701 16232
rect 5705 15763 8701 15796
rect 8849 15763 9629 16265
rect 9777 15763 10320 16265
rect 5705 15756 10320 15763
rect 840 15698 10320 15756
rect 400 15327 10322 15378
rect 400 15302 10113 15327
rect 400 15295 4753 15302
rect 400 14945 2797 15295
rect 3133 14950 4753 15295
rect 4945 14950 10113 15302
rect 3133 14946 10113 14950
rect 10259 14946 10322 15327
rect 3133 14945 10322 14946
rect 400 14877 10322 14945
rect 400 500 600 14877
rect 1193 14429 2349 14480
rect 1193 14250 1222 14429
rect 2301 14250 2349 14429
rect 1193 14207 2349 14250
rect 1663 650 1805 14207
rect 2390 13811 2596 13855
rect 2390 13290 2422 13811
rect 2562 13290 2596 13811
rect 2390 13241 2596 13290
rect 2441 1105 2546 13241
rect 2434 985 15271 1105
rect 1663 530 13339 650
rect 1663 529 1844 530
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 530
rect 15181 0 15271 985
use flashADC_3bit  flashADC_3bit_0
timestamp 1762640459
transform 1 0 2729 0 1 19824
box -1535 -5707 7777 2296
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel metal4 9139 22224 9169 22576 1 uo_out[1]
port 44 n
rlabel metal4 8863 22106 8893 22576 1 uo_out[2]
port 45 n
<< properties >>
string FIXED_BBOX 0 0 33488 22576
<< end >>
