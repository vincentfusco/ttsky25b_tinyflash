magic
tech sky130A
timestamp 1762723546
<< error_p >>
rect 10570 17920 10598 17934
rect 10584 17906 10598 17920
rect 4046 16968 4074 16982
rect 4060 16954 4074 16968
rect 4074 16912 4102 16926
rect 4088 16898 4102 16912
rect 4872 16898 4900 16912
rect 4872 16884 4914 16898
rect 4900 16870 4914 16884
rect 4844 16842 4872 16856
rect 4844 16828 4886 16842
rect 4872 16814 4886 16828
rect 4816 16786 4844 16800
rect 4130 16772 4158 16786
rect 4816 16772 4858 16786
rect 4144 16758 4158 16772
rect 4844 16758 4858 16772
rect 4788 16730 4816 16744
rect 4788 16716 4830 16730
rect 4816 16702 4830 16716
rect 4214 16632 4242 16646
rect 4228 16618 4242 16632
rect 4242 16576 4270 16590
rect 4256 16562 4270 16576
rect 4704 16534 4732 16548
rect 4270 16520 4298 16534
rect 4704 16520 4746 16534
rect 4284 16506 4298 16520
rect 4732 16506 4746 16520
rect 4676 16478 4704 16492
rect 4676 16464 4718 16478
rect 4704 16450 4718 16464
rect 4326 16436 4354 16450
rect 4340 16422 4354 16436
rect 4662 16408 4690 16422
rect 4676 16394 4690 16408
rect 4634 16352 4662 16366
rect 4648 16338 4662 16352
rect 3262 16212 3290 16226
rect 3262 16198 3276 16212
rect 4354 15316 4382 15330
rect 4354 15302 4368 15316
rect 4270 15260 4298 15274
rect 4270 15246 4284 15260
rect 4214 15232 4242 15246
rect 5838 15232 5866 15246
rect 4214 15218 4228 15232
rect 5852 15218 5866 15232
rect 4158 15204 4186 15218
rect 4158 15190 4172 15204
rect 3626 15176 3654 15190
rect 3640 15162 3654 15176
rect 4102 15176 4130 15190
rect 4102 15162 4116 15176
rect 4046 15148 4074 15162
rect 4046 15134 4060 15148
rect 3710 15092 3738 15106
rect 3724 15078 3738 15092
rect 3906 15092 3934 15106
rect 3906 15078 3920 15092
rect 9618 15064 9646 15078
rect 9632 15050 9646 15064
rect 9058 14840 9086 14854
rect 9058 14826 9072 14840
rect 9226 14700 9254 14714
rect 9240 14686 9254 14700
rect 9618 14672 9646 14686
rect 9618 14658 9632 14672
rect 9282 14616 9310 14630
rect 9296 14602 9310 14616
rect 9590 14616 9618 14630
rect 9590 14602 9604 14616
rect 9310 14588 9338 14602
rect 9324 14574 9338 14588
rect 9562 14588 9590 14602
rect 9562 14574 9576 14588
rect 4886 14560 4942 14574
rect 9338 14560 9366 14574
rect 4886 14546 4900 14560
rect 4928 14546 4942 14560
rect 9352 14546 9366 14560
rect 4746 14504 4774 14518
rect 4746 14490 4760 14504
rect 4690 14476 4718 14490
rect 4970 14476 4998 14490
rect 4690 14462 4704 14476
rect 4984 14462 4998 14476
rect 4634 14448 4662 14462
rect 4998 14448 5026 14462
rect 4634 14434 4648 14448
rect 5012 14434 5026 14448
rect 4578 14392 4606 14406
rect 4578 14378 4592 14392
rect 4970 14364 4998 14378
rect 9814 14364 9842 14378
rect 4970 14350 4984 14364
rect 9814 14350 9828 14364
rect 4914 14336 4942 14350
rect 9786 14336 9814 14350
rect 4914 14322 4928 14336
rect 9786 14322 9800 14336
rect 4858 14308 4886 14322
rect 4858 14294 4872 14308
rect 4802 14280 4830 14294
rect 9170 14280 9198 14294
rect 4802 14266 4816 14280
rect 9184 14266 9198 14280
rect 6762 14252 6790 14266
rect 10066 14252 10094 14266
rect 6762 14238 6776 14252
rect 10080 14238 10094 14252
rect 4662 14224 4690 14238
rect 6706 14224 6734 14238
rect 9086 14224 9114 14238
rect 4662 14210 4676 14224
rect 6706 14210 6720 14224
rect 9100 14210 9114 14224
rect 9590 14224 9618 14238
rect 9590 14210 9604 14224
rect 6818 14196 6846 14210
rect 6818 14182 6832 14196
rect 6818 14168 6846 14182
rect 6832 14154 6846 14168
rect 6006 14140 6034 14154
rect 6020 14126 6034 14140
rect 6818 14140 6846 14154
rect 7798 14140 7826 14154
rect 6818 14126 6832 14140
rect 7812 14126 7826 14140
rect 9534 14140 9562 14154
rect 9646 14140 9674 14154
rect 9534 14126 9548 14140
rect 9646 14126 9660 14140
rect 6034 14112 6062 14126
rect 6048 14098 6062 14112
rect 8582 14112 8610 14126
rect 9114 14112 9142 14126
rect 9198 14112 9226 14126
rect 8582 14098 8596 14112
rect 9128 14098 9142 14112
rect 9212 14098 9226 14112
rect 6874 14084 6902 14098
rect 6958 14084 7014 14098
rect 9506 14084 9534 14098
rect 9814 14084 9842 14098
rect 6874 14070 6888 14084
rect 6972 14070 7000 14084
rect 9506 14070 9520 14084
rect 9828 14070 9842 14084
rect 6874 14056 6902 14070
rect 6888 14042 6902 14056
rect 6958 14056 6986 14070
rect 9478 14056 9506 14070
rect 9590 14056 9618 14070
rect 6958 14042 6972 14056
rect 9478 14042 9492 14056
rect 9590 14042 9604 14056
rect 6874 14028 6902 14042
rect 8666 14028 8694 14042
rect 9842 14028 9870 14042
rect 6874 14014 6888 14028
rect 8680 14014 8694 14028
rect 9856 14014 9870 14028
rect 9142 14000 9170 14014
rect 9156 13986 9170 14000
rect 9450 14000 9478 14014
rect 9450 13986 9464 14000
rect 8302 13972 8330 13986
rect 8694 13972 8722 13986
rect 9226 13972 9254 13986
rect 8302 13958 8316 13972
rect 8708 13958 8722 13972
rect 9240 13958 9254 13972
rect 9534 13972 9562 13986
rect 9534 13958 9548 13972
rect 10066 13944 10094 13958
rect 10066 13930 10080 13944
rect 6174 13916 6202 13930
rect 8218 13916 8246 13930
rect 8722 13916 8750 13930
rect 6174 13902 6188 13916
rect 8218 13902 8232 13916
rect 8736 13902 8750 13916
rect 9114 13916 9142 13930
rect 9394 13916 9422 13930
rect 9506 13916 9534 13930
rect 9954 13916 9982 13930
rect 9114 13902 9128 13916
rect 9394 13902 9408 13916
rect 9506 13902 9520 13916
rect 9968 13902 9982 13916
rect 10038 13916 10066 13930
rect 10038 13902 10052 13916
rect 6118 13888 6146 13902
rect 8190 13888 8218 13902
rect 6118 13874 6132 13888
rect 8190 13874 8204 13888
rect 6678 13832 6706 13846
rect 6692 13818 6706 13832
rect 9338 13832 9366 13846
rect 9674 13832 9702 13846
rect 9338 13818 9352 13832
rect 9688 13818 9702 13832
rect 8134 13804 8162 13818
rect 9310 13804 9338 13818
rect 9506 13804 9534 13818
rect 9702 13804 9730 13818
rect 8134 13790 8148 13804
rect 9310 13790 9324 13804
rect 9506 13790 9520 13804
rect 9716 13790 9730 13804
rect 6706 13776 6734 13790
rect 6720 13762 6734 13776
rect 9478 13776 9506 13790
rect 9478 13762 9492 13776
rect 10122 13748 10150 13762
rect 10136 13734 10150 13748
rect 6734 13720 6762 13734
rect 6748 13706 6762 13720
rect 9450 13720 9478 13734
rect 10150 13720 10178 13734
rect 9450 13706 9464 13720
rect 10164 13706 10178 13720
rect 6482 13664 6510 13678
rect 6762 13664 6790 13678
rect 6482 13650 6496 13664
rect 6776 13650 6790 13664
rect 6426 13636 6454 13650
rect 6426 13622 6440 13636
rect 8134 13608 8162 13622
rect 9450 13608 9478 13622
rect 8148 13594 8162 13608
rect 9464 13594 9478 13608
rect 10150 13580 10178 13594
rect 10150 13566 10164 13580
rect 8162 13552 8190 13566
rect 8176 13538 8190 13552
rect 8498 13496 8526 13510
rect 9534 13496 9562 13510
rect 8498 13482 8512 13496
rect 9548 13482 9562 13496
rect 9646 13496 9674 13510
rect 9646 13482 9660 13496
rect 6622 13468 6650 13482
rect 6846 13468 6874 13482
rect 8246 13468 8274 13482
rect 6622 13454 6636 13468
rect 6860 13454 6874 13468
rect 8260 13454 8274 13468
rect 9562 13440 9590 13454
rect 9562 13426 9576 13440
rect 6874 13412 6902 13426
rect 6888 13398 6902 13412
rect 9562 13384 9590 13398
rect 9576 13370 9590 13384
rect 8218 13356 8246 13370
rect 8694 13356 8722 13370
rect 8218 13342 8232 13356
rect 8694 13342 8708 13356
rect 8638 13328 8666 13342
rect 9646 13328 9674 13342
rect 8638 13314 8652 13328
rect 9660 13314 9674 13328
rect 8218 13300 8246 13314
rect 8232 13286 8246 13300
rect 8582 13300 8610 13314
rect 9702 13300 9730 13314
rect 8582 13286 8596 13300
rect 9716 13286 9730 13300
rect 7798 13272 7826 13286
rect 8246 13272 8274 13286
rect 7798 13258 7812 13272
rect 8260 13258 8274 13272
rect 8526 13272 8554 13286
rect 8526 13258 8540 13272
rect 7770 13244 7798 13258
rect 9450 13244 9478 13258
rect 7770 13230 7784 13244
rect 9450 13230 9464 13244
rect 9422 13216 9450 13230
rect 9422 13202 9436 13216
rect 8302 13188 8330 13202
rect 8316 13174 8330 13188
rect 8582 13188 8610 13202
rect 8638 13188 8666 13202
rect 8582 13174 8596 13188
rect 8652 13174 8666 13188
rect 8330 13160 8358 13174
rect 8694 13160 8722 13174
rect 8344 13146 8358 13160
rect 8708 13146 8722 13160
rect 8722 13132 8750 13146
rect 9310 13132 9338 13146
rect 8736 13118 8750 13132
rect 9324 13118 9338 13132
rect 8778 13104 8806 13118
rect 9394 13104 9422 13118
rect 8792 13090 8806 13104
rect 9408 13090 9422 13104
rect 8806 13076 8834 13090
rect 9450 13076 9478 13090
rect 8820 13062 8834 13076
rect 9464 13062 9478 13076
rect 8834 13048 8862 13062
rect 8848 13034 8862 13048
rect 9282 13048 9310 13062
rect 9282 13034 9296 13048
rect 9590 13020 9618 13034
rect 9604 13006 9618 13020
rect 9646 13020 9674 13034
rect 9646 13006 9660 13020
rect 9142 12992 9170 13006
rect 9142 12978 9156 12992
rect 7994 12964 8022 12978
rect 8008 12950 8022 12964
rect 9086 12964 9114 12978
rect 9086 12950 9100 12964
rect 8302 12936 8330 12950
rect 8358 12936 8386 12950
rect 8302 12922 8316 12936
rect 8372 12922 8386 12936
rect 8778 12936 8806 12950
rect 8778 12922 8792 12936
rect 8274 12908 8302 12922
rect 8274 12894 8288 12908
rect 9030 12880 9058 12894
rect 9030 12866 9044 12880
rect 8050 12824 8078 12838
rect 8064 12810 8078 12824
rect 8190 12824 8218 12838
rect 8190 12810 8204 12824
rect 9002 12796 9030 12810
rect 9002 12782 9016 12796
rect 9366 12684 9394 12698
rect 9366 12670 9380 12684
rect 10178 12600 10206 12614
rect 10192 12586 10206 12600
rect 7742 12516 7770 12530
rect 10318 12516 10346 12530
rect 7756 12502 7770 12516
rect 10332 12502 10346 12516
rect 10402 12460 10430 12474
rect 10416 12446 10430 12460
rect 7770 12432 7798 12446
rect 7784 12418 7798 12432
rect 8022 12376 8050 12390
rect 8022 12362 8036 12376
rect 10626 12320 10654 12334
rect 10640 12306 10654 12320
rect 6650 12264 6678 12278
rect 6664 12250 6678 12264
rect 6286 12236 6314 12250
rect 6594 12236 6622 12250
rect 6300 12222 6314 12236
rect 6608 12222 6622 12236
rect 5922 12208 5950 12222
rect 6566 12208 6594 12222
rect 5936 12194 5950 12208
rect 6580 12194 6594 12208
rect 6258 12180 6286 12194
rect 6272 12166 6286 12180
rect 5950 12152 5978 12166
rect 6090 12152 6118 12166
rect 5964 12138 5978 12152
rect 6104 12138 6118 12152
rect 5922 12124 5950 12138
rect 5936 12110 5950 12124
rect 5726 12096 5754 12110
rect 5740 12082 5754 12096
rect 6174 12040 6202 12054
rect 6188 12026 6202 12040
rect 6034 11872 6062 11886
rect 6566 11872 6594 11886
rect 9142 11872 9170 11886
rect 6034 11858 6048 11872
rect 6566 11858 6580 11872
rect 9142 11858 9156 11872
rect 6482 11844 6510 11858
rect 9198 11844 9226 11858
rect 9506 11844 9534 11858
rect 6482 11830 6496 11844
rect 9198 11830 9212 11844
rect 9520 11830 9534 11844
rect 9226 11816 9254 11830
rect 9226 11802 9240 11816
rect 9254 11760 9282 11774
rect 9254 11746 9268 11760
rect 11634 11648 11662 11662
rect 11634 11634 11648 11648
rect 11662 11620 11690 11634
rect 13174 11620 13202 11634
rect 11662 11606 11676 11620
rect 13174 11606 13188 11620
rect 8274 11284 8302 11298
rect 8274 11270 8288 11284
rect 12810 11256 12838 11270
rect 12824 11242 12838 11256
rect 8078 11228 8106 11242
rect 8078 11214 8092 11228
rect 7994 11200 8022 11214
rect 7994 11186 8008 11200
rect 12838 11172 12866 11186
rect 12852 11158 12866 11172
rect 8218 11116 8246 11130
rect 8218 11102 8232 11116
rect 7994 11088 8022 11102
rect 8008 11074 8022 11088
rect 12838 11088 12894 11102
rect 12838 11074 12852 11088
rect 12880 11074 12894 11088
rect 8358 11032 8386 11046
rect 8372 11018 8386 11032
rect 8162 11004 8190 11018
rect 8176 10990 8190 11004
rect 12866 11004 12922 11018
rect 12866 10990 12880 11004
rect 12908 10990 12922 11004
rect 8022 10976 8050 10990
rect 8036 10962 8050 10976
rect 8386 10920 8414 10934
rect 8400 10906 8414 10920
rect 12894 10920 12950 10934
rect 12894 10906 12908 10920
rect 12936 10906 12950 10920
rect 8190 10892 8218 10906
rect 8204 10878 8218 10892
rect 8050 10864 8078 10878
rect 8064 10850 8078 10864
rect 10178 10836 10206 10850
rect 12950 10836 12978 10850
rect 10192 10822 10206 10836
rect 12964 10822 12978 10836
rect 8414 10808 8442 10822
rect 10066 10808 10094 10822
rect 8428 10794 8442 10808
rect 10080 10794 10094 10808
rect 8218 10780 8246 10794
rect 9954 10780 9982 10794
rect 8232 10766 8246 10780
rect 9968 10766 9982 10780
rect 8078 10752 8106 10766
rect 9842 10752 9870 10766
rect 12670 10752 12698 10766
rect 8092 10738 8106 10752
rect 9856 10738 9870 10752
rect 12684 10738 12698 10752
rect 9730 10724 9758 10738
rect 9744 10710 9758 10724
rect 12558 10724 12586 10738
rect 12558 10710 12572 10724
rect 8442 10696 8470 10710
rect 9618 10696 9646 10710
rect 8456 10682 8470 10696
rect 9632 10682 9646 10696
rect 8246 10668 8274 10682
rect 9506 10668 9534 10682
rect 8260 10654 8274 10668
rect 9520 10654 9534 10668
rect 12726 10668 12754 10682
rect 12726 10654 12740 10668
rect 9394 10640 9422 10654
rect 9408 10626 9422 10640
rect 10346 10640 10374 10654
rect 12838 10640 12866 10654
rect 10346 10626 10360 10640
rect 12852 10626 12866 10640
rect 12418 10612 12446 10626
rect 12432 10598 12446 10612
rect 12474 10612 12502 10626
rect 12474 10598 12488 10612
rect 8470 10584 8498 10598
rect 8484 10570 8498 10584
rect 12642 10584 12670 10598
rect 12642 10570 12656 10584
rect 8134 10556 8162 10570
rect 8274 10556 8302 10570
rect 8148 10542 8162 10556
rect 8288 10542 8302 10556
rect 12614 10556 12642 10570
rect 12614 10542 12628 10556
rect 10374 10528 10402 10542
rect 10374 10514 10388 10528
rect 12390 10500 12418 10514
rect 12390 10486 12404 10500
rect 8498 10472 8526 10486
rect 8512 10458 8526 10472
rect 12362 10472 12390 10486
rect 12362 10458 12376 10472
rect 8162 10444 8190 10458
rect 8302 10444 8330 10458
rect 8176 10430 8190 10444
rect 8316 10430 8330 10444
rect 8526 10360 8554 10374
rect 8540 10346 8554 10360
rect 8190 10332 8218 10346
rect 8330 10332 8358 10346
rect 8204 10318 8218 10332
rect 8344 10318 8358 10332
rect 10766 10276 10794 10290
rect 10780 10262 10794 10276
rect 8554 10248 8582 10262
rect 9114 10248 9142 10262
rect 8568 10234 8582 10248
rect 9128 10234 9142 10248
rect 8218 10220 8246 10234
rect 9366 10220 9394 10234
rect 8232 10206 8246 10220
rect 9380 10206 9394 10220
rect 10038 10192 10066 10206
rect 10052 10178 10066 10192
rect 11494 10192 11522 10206
rect 11494 10178 11508 10192
rect 8386 10136 8414 10150
rect 8400 10122 8414 10136
rect 8470 10136 8498 10150
rect 9114 10136 9142 10150
rect 9618 10136 9646 10150
rect 9954 10136 9982 10150
rect 8470 10122 8484 10136
rect 9114 10122 9128 10136
rect 9618 10122 9632 10136
rect 9954 10122 9968 10136
rect 8246 10108 8274 10122
rect 8260 10094 8274 10108
rect 9842 10108 9870 10122
rect 9842 10094 9856 10108
rect 9562 10080 9618 10094
rect 9562 10066 9576 10080
rect 9604 10066 9618 10080
rect 9702 10080 9730 10094
rect 10038 10080 10066 10094
rect 12418 10080 12446 10094
rect 9702 10066 9716 10080
rect 10038 10066 10052 10080
rect 12432 10066 12446 10080
rect 8666 10052 8694 10066
rect 9590 10052 9618 10066
rect 9926 10052 9954 10066
rect 10150 10052 10178 10066
rect 8666 10038 8680 10052
rect 9590 10038 9604 10052
rect 9926 10038 9940 10052
rect 10164 10038 10178 10052
rect 8274 10024 8302 10038
rect 8288 10010 8302 10024
rect 8638 10024 8666 10038
rect 9786 10024 9814 10038
rect 8638 10010 8652 10024
rect 9786 10010 9800 10024
rect 8610 9996 8638 10010
rect 9674 9996 9702 10010
rect 8610 9982 8624 9996
rect 9674 9982 9688 9996
rect 9562 9968 9590 9982
rect 9562 9954 9576 9968
rect 10822 9940 10850 9954
rect 10822 9926 10836 9940
rect 10318 9912 10346 9926
rect 10332 9898 10346 9912
rect 10990 9884 11018 9898
rect 10990 9870 11004 9884
rect 11942 9828 11970 9842
rect 11956 9814 11970 9828
rect 13454 9772 13482 9786
rect 13874 9772 13902 9786
rect 13454 9758 13468 9772
rect 13888 9758 13902 9772
rect 9226 9744 9254 9758
rect 12138 9744 12166 9758
rect 9240 9730 9254 9744
rect 12152 9730 12166 9744
rect 13370 9744 13398 9758
rect 13370 9730 13384 9744
rect 10178 9716 10206 9730
rect 13314 9716 13342 9730
rect 13762 9716 13790 9730
rect 10178 9702 10192 9716
rect 13314 9702 13328 9716
rect 13762 9702 13776 9716
rect 9562 9688 9590 9702
rect 9576 9674 9590 9688
rect 10150 9688 10178 9702
rect 10150 9674 10164 9688
rect 9590 9632 9618 9646
rect 12698 9632 12726 9646
rect 9604 9618 9618 9632
rect 12712 9618 12726 9632
rect 9618 9604 9646 9618
rect 12754 9604 12782 9618
rect 9632 9590 9646 9604
rect 12768 9590 12782 9604
rect 7126 9352 7154 9366
rect 7140 9338 7154 9352
rect 7070 9324 7098 9338
rect 7084 9310 7098 9324
rect 7014 9296 7042 9310
rect 7028 9282 7042 9296
rect 6958 9268 6986 9282
rect 6972 9254 6986 9268
rect 6902 9240 6930 9254
rect 6916 9226 6930 9240
rect 5782 9212 5810 9226
rect 9394 9212 9422 9226
rect 5782 9198 5796 9212
rect 9408 9198 9422 9212
rect 12194 9100 12222 9114
rect 12208 9086 12222 9100
rect 5586 9072 5614 9086
rect 9450 9072 9478 9086
rect 5586 9058 5600 9072
rect 9464 9058 9478 9072
rect 12166 9044 12194 9058
rect 12180 9030 12194 9044
rect 9478 9016 9506 9030
rect 9492 9002 9506 9016
rect 9534 8988 9562 9002
rect 12138 8988 12166 9002
rect 9534 8974 9548 8988
rect 12152 8974 12166 8988
rect 9534 8932 9562 8946
rect 12110 8932 12138 8946
rect 9548 8918 9562 8932
rect 12124 8904 12152 8932
rect 12082 8876 12110 8890
rect 12096 8848 12124 8876
rect 12054 8820 12082 8834
rect 12068 8792 12096 8820
rect 12026 8764 12054 8778
rect 5530 8736 5558 8750
rect 12040 8736 12068 8764
rect 5544 8722 5558 8736
rect 11606 8708 11634 8722
rect 11998 8708 12026 8722
rect 11620 8694 11634 8708
rect 12012 8694 12026 8708
rect 5558 8680 5586 8694
rect 11326 8680 11354 8694
rect 5572 8666 5586 8680
rect 11340 8666 11354 8680
rect 11970 8652 11998 8666
rect 11984 8638 11998 8652
rect 6202 8624 6230 8638
rect 6202 8610 6216 8624
rect 11942 8596 11970 8610
rect 11956 8582 11970 8596
rect 5642 8568 5670 8582
rect 5656 8554 5670 8568
rect 6062 8512 6090 8526
rect 6062 8498 6076 8512
rect 6006 8484 6034 8498
rect 6006 8470 6020 8484
rect 6510 8120 6538 8134
rect 6510 8106 6524 8120
rect 6538 8092 6566 8106
rect 6538 8078 6552 8092
rect 5362 8064 5390 8078
rect 5376 8050 5390 8064
rect 6594 8008 6622 8022
rect 6594 7994 6608 8008
rect 5306 7980 5334 7994
rect 5320 7966 5334 7980
rect 6622 7980 6650 7994
rect 6622 7966 6636 7980
rect 5250 7896 5278 7910
rect 5264 7882 5278 7896
rect 6678 7896 6706 7910
rect 6678 7882 6692 7896
rect 6706 7868 6734 7882
rect 6706 7854 6720 7868
rect 5194 7812 5222 7826
rect 5208 7798 5222 7812
rect 6734 7812 6762 7826
rect 6734 7798 6748 7812
rect 5166 7784 5194 7798
rect 5180 7770 5194 7784
rect 5138 7728 5166 7742
rect 5152 7714 5166 7728
rect 10934 6104 10962 6118
rect 10948 6090 10962 6104
rect 9786 5544 9814 5558
rect 9786 5530 9800 5544
rect 13790 5348 13818 5362
rect 13804 5334 13818 5348
rect 13650 5320 13678 5334
rect 13846 5320 13874 5334
rect 13650 5306 13664 5320
rect 13860 5306 13874 5320
rect 13986 5264 14014 5278
rect 14000 5250 14014 5264
rect 14042 5236 14070 5250
rect 14056 5222 14070 5236
rect 14098 5208 14126 5222
rect 14112 5194 14126 5208
rect 14154 5180 14182 5194
rect 14168 5166 14182 5180
rect 14238 5152 14266 5166
rect 14252 5138 14266 5152
rect 14238 5124 14266 5138
rect 14322 5152 14350 5166
rect 14322 5138 14336 5152
rect 14322 5124 14350 5138
rect 14238 5110 14252 5124
rect 14336 5110 14350 5124
rect 14714 5068 14742 5082
rect 14728 5054 14742 5068
rect 14770 5040 14798 5054
rect 14784 5026 14798 5040
rect 14798 5012 14826 5026
rect 14812 4998 14826 5012
rect 14826 4984 14854 4998
rect 14840 4970 14854 4984
<< metal2 >>
rect 6944 17920 7224 17948
rect 6944 17892 7252 17920
rect 6944 17864 7280 17892
rect 6944 17836 7028 17864
rect 7168 17836 7280 17864
rect 7392 17836 7476 17948
rect 7840 17892 7980 17948
rect 7812 17864 7980 17892
rect 7812 17836 7868 17864
rect 6916 17808 7028 17836
rect 3668 17724 3836 17752
rect 3584 17696 3836 17724
rect 6916 17696 7000 17808
rect 7196 17780 7280 17836
rect 7364 17808 7476 17836
rect 3528 17668 3836 17696
rect 3500 17640 3836 17668
rect 3472 17556 3808 17640
rect 6888 17584 6972 17696
rect 7168 17640 7252 17780
rect 7364 17696 7448 17808
rect 7784 17752 7868 17836
rect 7140 17612 7224 17640
rect 7112 17584 7224 17612
rect 4396 17556 4592 17584
rect 6888 17556 7196 17584
rect 7336 17556 7420 17696
rect 7756 17668 7840 17752
rect 7728 17612 7812 17668
rect 7896 17612 7980 17864
rect 8176 17836 8260 17948
rect 8456 17920 8568 17948
rect 8624 17920 8904 17948
rect 8456 17892 8540 17920
rect 8428 17864 8512 17892
rect 8148 17808 8260 17836
rect 8400 17836 8512 17864
rect 8624 17864 8876 17920
rect 8624 17836 8708 17864
rect 9184 17836 9352 17948
rect 9548 17892 9716 17948
rect 9912 17920 10108 17948
rect 10276 17920 10584 17948
rect 10612 17920 10920 17948
rect 9884 17892 10136 17920
rect 8400 17808 8484 17836
rect 8596 17808 8708 17836
rect 8148 17696 8232 17808
rect 8372 17752 8456 17808
rect 8344 17724 8428 17752
rect 8316 17696 8428 17724
rect 8596 17696 8680 17808
rect 9156 17696 9240 17836
rect 9296 17808 9352 17836
rect 9520 17836 9716 17892
rect 9828 17864 10136 17892
rect 10248 17864 10556 17920
rect 10584 17864 10892 17920
rect 9828 17836 9940 17864
rect 9520 17808 9576 17836
rect 7728 17584 7784 17612
rect 7896 17584 7952 17612
rect 3444 17332 3808 17556
rect 4340 17528 4424 17556
rect 4312 17500 4368 17528
rect 4564 17500 4592 17556
rect 4256 17472 4340 17500
rect 4536 17472 4592 17500
rect 6860 17500 7168 17556
rect 4228 17444 4284 17472
rect 4508 17444 4564 17472
rect 6860 17444 6944 17500
rect 7084 17472 7196 17500
rect 4172 17416 4256 17444
rect 4480 17416 4536 17444
rect 6832 17416 6944 17444
rect 7112 17444 7224 17472
rect 7308 17444 7392 17556
rect 7700 17528 7784 17584
rect 7672 17444 7756 17528
rect 4144 17388 4200 17416
rect 4452 17388 4508 17416
rect 4116 17360 4172 17388
rect 4396 17360 4480 17388
rect 4060 17332 4144 17360
rect 4368 17332 4452 17360
rect 3416 17304 3808 17332
rect 4032 17304 4088 17332
rect 4340 17304 4396 17332
rect 6832 17304 6916 17416
rect 7112 17332 7196 17444
rect 7280 17416 7392 17444
rect 7644 17416 7728 17444
rect 7868 17416 7952 17584
rect 8120 17584 8204 17696
rect 8316 17668 8400 17696
rect 8288 17612 8372 17668
rect 8260 17584 8344 17612
rect 8568 17584 8652 17696
rect 8120 17556 8316 17584
rect 8568 17556 8792 17584
rect 9128 17556 9212 17696
rect 9268 17668 9352 17808
rect 9492 17752 9576 17808
rect 9492 17724 9548 17752
rect 9604 17724 9688 17836
rect 9800 17808 9912 17836
rect 9800 17724 9884 17808
rect 9464 17668 9548 17724
rect 8092 17500 8316 17556
rect 8092 17444 8176 17500
rect 3416 17192 3780 17304
rect 4004 17276 4060 17304
rect 4312 17276 4368 17304
rect 3976 17248 4032 17276
rect 4284 17248 4340 17276
rect 3948 17220 4004 17248
rect 4256 17220 4312 17248
rect 3892 17192 3976 17220
rect 4228 17192 4284 17220
rect 3416 17164 3724 17192
rect 3864 17164 3920 17192
rect 4200 17164 4256 17192
rect 4844 17164 5236 17248
rect 6804 17192 6888 17304
rect 7084 17220 7168 17332
rect 7280 17304 7364 17416
rect 7644 17360 7952 17416
rect 7616 17332 7952 17360
rect 7028 17192 7168 17220
rect 7252 17192 7336 17304
rect 7616 17276 7700 17332
rect 7588 17220 7672 17276
rect 7560 17192 7672 17220
rect 7868 17192 7952 17332
rect 8064 17416 8176 17444
rect 8232 17444 8316 17500
rect 8540 17500 8792 17556
rect 8540 17444 8624 17500
rect 9100 17444 9184 17556
rect 9268 17500 9324 17668
rect 9464 17640 9520 17668
rect 9436 17584 9520 17640
rect 9576 17584 9660 17724
rect 9772 17696 9884 17724
rect 10052 17780 10164 17864
rect 10360 17780 10444 17864
rect 10696 17780 10780 17864
rect 9772 17584 9856 17696
rect 10052 17668 10136 17780
rect 10332 17668 10416 17780
rect 10668 17668 10752 17780
rect 9436 17556 9492 17584
rect 8064 17304 8148 17416
rect 8232 17388 8344 17444
rect 8260 17304 8344 17388
rect 8512 17416 8624 17444
rect 9072 17416 9184 17444
rect 8512 17304 8596 17416
rect 9072 17304 9156 17416
rect 9240 17360 9324 17500
rect 9408 17500 9492 17556
rect 9408 17472 9464 17500
rect 9548 17472 9632 17584
rect 9380 17416 9464 17472
rect 9520 17444 9632 17472
rect 9744 17444 9828 17584
rect 10024 17528 10108 17668
rect 10304 17640 10416 17668
rect 10640 17640 10752 17668
rect 10304 17528 10388 17640
rect 10640 17528 10724 17640
rect 9380 17388 9436 17416
rect 6804 17164 7140 17192
rect 7252 17164 7504 17192
rect 3416 17136 3668 17164
rect 3836 17136 3892 17164
rect 4144 17136 4228 17164
rect 3388 17108 3612 17136
rect 3808 17108 3864 17136
rect 4116 17108 4200 17136
rect 3388 17052 3556 17108
rect 3780 17080 3836 17108
rect 4088 17080 4172 17108
rect 3752 17052 3808 17080
rect 4060 17052 4144 17080
rect 3388 17024 3528 17052
rect 3724 17024 3780 17052
rect 4032 17024 4116 17052
rect 3360 16996 3528 17024
rect 3696 16996 3752 17024
rect 4004 16996 4060 17024
rect 4844 16996 4900 17164
rect 3360 16968 3500 16996
rect 3668 16968 3724 16996
rect 3976 16968 4060 16996
rect 3332 16912 3500 16968
rect 3640 16940 3696 16968
rect 3948 16940 4004 16968
rect 3612 16912 3668 16940
rect 3920 16912 3976 16940
rect 4060 16912 4088 16968
rect 4816 16912 4900 16996
rect 3332 16828 3472 16912
rect 3584 16884 3640 16912
rect 3864 16884 3948 16912
rect 3556 16856 3612 16884
rect 3836 16856 3920 16884
rect 4088 16856 4116 16912
rect 4788 16884 4900 16912
rect 4928 17080 5236 17164
rect 6776 17136 7112 17164
rect 6776 17108 7056 17136
rect 7224 17108 7476 17164
rect 7560 17136 7644 17192
rect 7840 17136 7952 17192
rect 8036 17164 8120 17304
rect 8260 17248 8372 17304
rect 8288 17164 8372 17248
rect 8484 17192 8568 17304
rect 8484 17164 8736 17192
rect 9044 17164 9128 17304
rect 9240 17192 9296 17360
rect 9352 17332 9436 17388
rect 9520 17332 9604 17444
rect 9716 17332 9800 17444
rect 9996 17416 10080 17528
rect 9352 17304 9408 17332
rect 9324 17248 9408 17304
rect 9324 17192 9380 17248
rect 9492 17192 9576 17332
rect 9688 17304 9800 17332
rect 9968 17388 10080 17416
rect 10276 17500 10388 17528
rect 10612 17500 10724 17528
rect 10276 17388 10360 17500
rect 10612 17388 10696 17500
rect 9688 17220 9772 17304
rect 9968 17276 10052 17388
rect 9940 17248 10052 17276
rect 10248 17248 10332 17388
rect 10584 17248 10668 17388
rect 9940 17220 10024 17248
rect 9688 17192 9800 17220
rect 9912 17192 10024 17220
rect 9212 17164 9380 17192
rect 7532 17108 7616 17136
rect 7840 17108 7924 17136
rect 8008 17108 8092 17164
rect 8288 17108 8400 17164
rect 8456 17108 8736 17164
rect 9016 17108 9100 17164
rect 9212 17108 9352 17164
rect 9464 17108 9548 17192
rect 9688 17164 9996 17192
rect 9716 17136 9968 17164
rect 10220 17136 10304 17248
rect 10556 17136 10640 17248
rect 9744 17108 9940 17136
rect 10192 17108 10304 17136
rect 10528 17108 10640 17136
rect 4928 17052 5264 17080
rect 4928 17024 5488 17052
rect 4928 16996 5544 17024
rect 4928 16968 5628 16996
rect 4928 16940 5684 16968
rect 4928 16912 5740 16940
rect 4928 16884 5796 16912
rect 4788 16856 4872 16884
rect 3528 16828 3584 16856
rect 3808 16828 3892 16856
rect 4088 16828 4144 16856
rect 3304 16800 3556 16828
rect 3780 16800 3864 16828
rect 3304 16716 3528 16800
rect 3724 16772 3836 16800
rect 4116 16772 4144 16828
rect 4760 16828 4872 16856
rect 4900 16856 5852 16884
rect 6720 16856 10696 16940
rect 4900 16828 5908 16856
rect 4760 16800 4844 16828
rect 4732 16772 4844 16800
rect 4872 16800 5992 16828
rect 6692 16800 10668 16856
rect 4872 16772 6048 16800
rect 3696 16744 3808 16772
rect 3612 16716 3808 16744
rect 4144 16744 4172 16772
rect 4732 16744 4816 16772
rect 4144 16716 4200 16744
rect 3304 16688 3696 16716
rect 3304 16660 3640 16688
rect 3752 16660 3808 16716
rect 4172 16688 4200 16716
rect 4704 16716 4816 16744
rect 4844 16744 6104 16772
rect 6692 16744 10640 16800
rect 4844 16716 5376 16744
rect 5488 16716 6160 16744
rect 6692 16716 10612 16744
rect 4704 16688 4788 16716
rect 4172 16660 4228 16688
rect 3332 16604 3668 16660
rect 3752 16604 3836 16660
rect 4200 16632 4228 16660
rect 4676 16660 4788 16688
rect 4816 16660 5348 16716
rect 5572 16688 6160 16716
rect 5684 16660 6160 16688
rect 4676 16632 5320 16660
rect 5796 16632 6160 16660
rect 3304 16576 3640 16604
rect 3780 16576 3864 16604
rect 4228 16576 4256 16632
rect 4648 16604 4760 16632
rect 4788 16604 5320 16632
rect 5880 16604 6132 16632
rect 4648 16576 5320 16604
rect 3276 16520 3640 16576
rect 3808 16548 3892 16576
rect 3248 16492 3304 16520
rect 3332 16492 3640 16520
rect 3836 16520 3920 16548
rect 4256 16520 4284 16576
rect 4620 16520 4732 16576
rect 4760 16520 5292 16576
rect 3836 16492 3976 16520
rect 4284 16492 4312 16520
rect 3220 16464 3276 16492
rect 3332 16464 3612 16492
rect 3892 16464 4032 16492
rect 4284 16464 4340 16492
rect 4592 16464 4704 16520
rect 4732 16464 5320 16520
rect 3192 16408 3248 16464
rect 3360 16436 3612 16464
rect 3920 16436 4116 16464
rect 4312 16436 4340 16464
rect 3360 16408 3584 16436
rect 3976 16408 4228 16436
rect 4340 16408 4368 16436
rect 4564 16408 4676 16464
rect 4704 16408 5348 16464
rect 6216 16436 6888 16464
rect 5880 16408 7588 16436
rect 3164 16380 3220 16408
rect 3360 16380 3556 16408
rect 4060 16380 4396 16408
rect 3136 16324 3192 16380
rect 3360 16352 3528 16380
rect 4144 16352 4424 16380
rect 4536 16352 4648 16408
rect 4676 16352 5348 16408
rect 5796 16380 7868 16408
rect 5740 16352 5964 16380
rect 7476 16352 8008 16380
rect 3388 16324 3500 16352
rect 4256 16324 4620 16352
rect 4648 16324 5348 16352
rect 5684 16324 5852 16352
rect 7812 16324 8064 16352
rect 3108 16268 3164 16324
rect 4340 16296 5348 16324
rect 5656 16296 5768 16324
rect 7980 16296 8092 16324
rect 3304 16268 3332 16296
rect 4424 16268 5320 16296
rect 5628 16268 5740 16296
rect 8036 16268 8120 16296
rect 3080 16212 3136 16268
rect 3276 16240 3332 16268
rect 4508 16240 5320 16268
rect 5600 16240 5684 16268
rect 8064 16240 8148 16268
rect 3276 16212 3304 16240
rect 3892 16212 3920 16240
rect 4592 16212 5320 16240
rect 5572 16212 5656 16240
rect 8092 16212 8176 16240
rect 3052 16156 3108 16212
rect 3248 16184 3276 16212
rect 3836 16184 3920 16212
rect 4676 16184 5292 16212
rect 5544 16184 5628 16212
rect 3220 16156 3276 16184
rect 3808 16156 3892 16184
rect 4732 16156 5292 16184
rect 5516 16156 5600 16184
rect 7644 16156 7980 16184
rect 8120 16156 8204 16212
rect 3024 16100 3080 16156
rect 3220 16128 3248 16156
rect 3752 16128 3864 16156
rect 4816 16128 5292 16156
rect 2996 16072 3080 16100
rect 3192 16100 3248 16128
rect 3724 16100 3808 16128
rect 4900 16100 5292 16128
rect 5488 16100 5572 16156
rect 6580 16128 6972 16156
rect 7476 16128 8064 16156
rect 8148 16128 8232 16156
rect 6384 16100 6664 16128
rect 7336 16100 7644 16128
rect 7924 16100 8092 16128
rect 8176 16100 8260 16128
rect 3192 16072 3220 16100
rect 3696 16072 3780 16100
rect 4984 16072 5264 16100
rect 5460 16072 5544 16100
rect 6244 16072 6496 16100
rect 7224 16072 7476 16100
rect 8008 16072 8120 16100
rect 8204 16072 8288 16100
rect 2996 16016 3052 16072
rect 3164 16044 3220 16072
rect 3640 16044 3752 16072
rect 5068 16044 5348 16072
rect 5460 16044 5516 16072
rect 6104 16044 6356 16072
rect 7112 16044 7336 16072
rect 8036 16044 8120 16072
rect 8232 16044 8316 16072
rect 3164 16016 3192 16044
rect 3612 16016 3696 16044
rect 5180 16016 5516 16044
rect 5992 16016 6244 16044
rect 7028 16016 7196 16044
rect 8064 16016 8120 16044
rect 8260 16016 8316 16044
rect 2968 15932 3024 16016
rect 3136 15988 3192 16016
rect 3584 15988 3668 16016
rect 5264 15988 5600 16016
rect 5880 15988 6132 16016
rect 6944 15988 7084 16016
rect 3136 15960 3164 15988
rect 3556 15960 3640 15988
rect 5376 15960 6020 15988
rect 6860 15960 7000 15988
rect 2940 15904 3024 15932
rect 3108 15904 3164 15960
rect 3528 15932 3612 15960
rect 5516 15932 5908 15960
rect 6776 15932 6916 15960
rect 8064 15932 8148 16016
rect 8260 15988 8344 16016
rect 8288 15960 8372 15988
rect 8316 15932 8400 15960
rect 3500 15904 3584 15932
rect 5488 15904 5712 15932
rect 5768 15904 5880 15932
rect 6720 15904 6832 15932
rect 8092 15904 8176 15932
rect 8344 15904 8400 15932
rect 2940 15820 2996 15904
rect 3108 15876 3136 15904
rect 3472 15876 3556 15904
rect 5404 15876 5628 15904
rect 5796 15876 5908 15904
rect 6636 15876 6748 15904
rect 8092 15876 8204 15904
rect 8344 15876 8428 15904
rect 3080 15820 3136 15876
rect 3444 15848 3528 15876
rect 5292 15848 5544 15876
rect 5824 15848 5936 15876
rect 6580 15848 6664 15876
rect 8120 15848 8204 15876
rect 8372 15848 8456 15876
rect 3416 15820 3500 15848
rect 5208 15820 5432 15848
rect 5852 15820 5964 15848
rect 6580 15820 6608 15848
rect 8120 15820 8232 15848
rect 8400 15820 8484 15848
rect 2912 15792 2996 15820
rect 2912 15652 2968 15792
rect 3052 15736 3108 15820
rect 3416 15792 3472 15820
rect 5124 15792 5348 15820
rect 5908 15792 5992 15820
rect 8148 15792 8260 15820
rect 8428 15792 8484 15820
rect 3388 15764 3444 15792
rect 5040 15764 5264 15792
rect 5936 15764 6048 15792
rect 8176 15764 8288 15792
rect 8428 15764 8512 15792
rect 3360 15736 3444 15764
rect 4956 15736 5180 15764
rect 5964 15736 6076 15764
rect 8204 15736 8344 15764
rect 8456 15736 8540 15764
rect 3052 15708 3080 15736
rect 2884 15540 2968 15652
rect 3024 15596 3080 15708
rect 3332 15708 3416 15736
rect 4872 15708 5068 15736
rect 5992 15708 6104 15736
rect 8232 15708 8372 15736
rect 8428 15708 8540 15736
rect 3332 15680 3388 15708
rect 4760 15680 4984 15708
rect 6020 15680 6160 15708
rect 8260 15680 8568 15708
rect 3304 15652 3388 15680
rect 4676 15652 4900 15680
rect 6076 15652 6216 15680
rect 8288 15652 8484 15680
rect 8512 15652 8596 15680
rect 3304 15624 3360 15652
rect 4592 15624 4816 15652
rect 6104 15624 6272 15652
rect 8288 15624 8428 15652
rect 8540 15624 8624 15652
rect 3276 15596 3332 15624
rect 4508 15596 4732 15624
rect 6160 15596 6328 15624
rect 8232 15596 8372 15624
rect 8568 15596 8624 15624
rect 2884 15372 2940 15540
rect 2884 15288 2968 15372
rect 2996 15288 3052 15596
rect 3248 15568 3332 15596
rect 4424 15568 4648 15596
rect 5684 15568 5740 15596
rect 6216 15568 6356 15596
rect 8204 15568 8344 15596
rect 8596 15568 8652 15596
rect 3248 15540 3304 15568
rect 4340 15540 4564 15568
rect 5628 15540 5712 15568
rect 6272 15540 6356 15568
rect 8176 15540 8288 15568
rect 8596 15540 8680 15568
rect 3220 15512 3304 15540
rect 4256 15512 4480 15540
rect 5544 15512 5656 15540
rect 6300 15512 6356 15540
rect 8120 15512 8260 15540
rect 8624 15512 8680 15540
rect 3220 15456 3276 15512
rect 4172 15484 4396 15512
rect 5488 15484 5600 15512
rect 4088 15456 4284 15484
rect 3192 15400 3248 15456
rect 4004 15428 4200 15456
rect 3920 15400 4116 15428
rect 3164 15372 3248 15400
rect 3836 15372 4032 15400
rect 3164 15316 3220 15372
rect 3752 15344 3948 15372
rect 3668 15316 3864 15344
rect 4368 15316 4396 15484
rect 5404 15456 5544 15484
rect 6132 15456 6188 15484
rect 6300 15456 6384 15512
rect 8092 15484 8204 15512
rect 8652 15484 8708 15512
rect 8064 15456 8176 15484
rect 5348 15428 5460 15456
rect 6076 15428 6160 15456
rect 5264 15400 5404 15428
rect 6020 15400 6132 15428
rect 5208 15372 5348 15400
rect 5964 15372 6104 15400
rect 6328 15372 6384 15456
rect 8036 15428 8148 15456
rect 8680 15428 8736 15484
rect 8008 15400 8120 15428
rect 8708 15400 8764 15428
rect 5124 15344 5292 15372
rect 5908 15344 6076 15372
rect 5068 15316 5236 15344
rect 5880 15316 6048 15344
rect 2884 15232 3052 15288
rect 3136 15288 3220 15316
rect 3584 15288 3780 15316
rect 4312 15288 4368 15316
rect 4984 15288 5180 15316
rect 5824 15288 6020 15316
rect 2912 15204 3080 15232
rect 3136 15204 3192 15288
rect 3500 15260 3696 15288
rect 4284 15260 4340 15288
rect 4928 15260 5124 15288
rect 5768 15260 5992 15288
rect 3416 15232 3612 15260
rect 4228 15232 4284 15260
rect 4844 15232 5068 15260
rect 5712 15232 5852 15260
rect 5880 15232 5964 15260
rect 6328 15232 6412 15372
rect 8008 15344 8092 15400
rect 8736 15372 8792 15400
rect 8036 15288 8120 15344
rect 8764 15316 8820 15372
rect 8792 15288 8848 15316
rect 8064 15260 8148 15288
rect 8820 15260 8876 15288
rect 8092 15232 8176 15260
rect 3332 15204 3528 15232
rect 3584 15204 3640 15232
rect 4172 15204 4228 15232
rect 4788 15204 4984 15232
rect 5656 15204 5796 15232
rect 5852 15204 5936 15232
rect 2968 15176 3192 15204
rect 3248 15176 3444 15204
rect 3612 15176 3640 15204
rect 4116 15176 4172 15204
rect 4732 15176 4928 15204
rect 5600 15176 5740 15204
rect 5824 15176 5908 15204
rect 6328 15176 6384 15232
rect 8120 15204 8204 15232
rect 8148 15176 8232 15204
rect 9520 15176 9576 15204
rect 2996 15148 3388 15176
rect 3640 15148 3668 15176
rect 4060 15148 4116 15176
rect 4648 15148 4872 15176
rect 5544 15148 5684 15176
rect 5796 15148 5880 15176
rect 6300 15148 6412 15176
rect 8176 15148 8260 15176
rect 9492 15148 9604 15176
rect 3052 15120 3304 15148
rect 3640 15120 3696 15148
rect 3976 15120 4060 15148
rect 4592 15120 4816 15148
rect 5488 15120 5628 15148
rect 5796 15120 5852 15148
rect 6272 15120 6440 15148
rect 8204 15120 8288 15148
rect 9464 15120 9632 15148
rect 3080 15092 3248 15120
rect 3668 15092 3724 15120
rect 3920 15092 4004 15120
rect 4508 15092 4760 15120
rect 5460 15092 5572 15120
rect 5768 15092 5824 15120
rect 6272 15092 6356 15120
rect 6412 15092 6496 15120
rect 8232 15092 8316 15120
rect 9408 15092 9576 15120
rect 3108 15064 3304 15092
rect 3724 15064 3920 15092
rect 4452 15064 4704 15092
rect 5404 15064 5516 15092
rect 5740 15064 5796 15092
rect 6272 15064 6328 15092
rect 6468 15064 6524 15092
rect 8176 15064 8344 15092
rect 9380 15064 9548 15092
rect 9604 15064 9632 15120
rect 3164 15036 3332 15064
rect 4368 15036 4648 15064
rect 5348 15036 5460 15064
rect 5712 15036 5768 15064
rect 3220 15008 3360 15036
rect 4312 15008 4592 15036
rect 5292 15008 5404 15036
rect 5684 15008 5740 15036
rect 3248 14980 3416 15008
rect 4228 14980 4508 15008
rect 5236 14980 5348 15008
rect 5656 14980 5712 15008
rect 6244 14980 6328 15064
rect 6496 15036 6580 15064
rect 8120 15036 8232 15064
rect 8288 15036 8372 15064
rect 9352 15036 9520 15064
rect 6524 15008 6608 15036
rect 8036 15008 8148 15036
rect 8316 15008 8400 15036
rect 9324 15008 9492 15036
rect 6580 14980 6636 15008
rect 7952 14980 8092 15008
rect 8344 14980 8428 15008
rect 9296 14980 9464 15008
rect 3276 14952 3444 14980
rect 4172 14952 4452 14980
rect 5180 14952 5292 14980
rect 5628 14952 5712 14980
rect 6272 14952 6328 14980
rect 6608 14952 6692 14980
rect 7868 14952 8008 14980
rect 8400 14952 8456 14980
rect 9268 14952 9436 14980
rect 3332 14924 3500 14952
rect 4088 14924 4396 14952
rect 5124 14924 5236 14952
rect 5628 14924 5684 14952
rect 6272 14924 6356 14952
rect 6664 14924 6720 14952
rect 7812 14924 7924 14952
rect 8428 14924 8484 14952
rect 9240 14924 9408 14952
rect 9632 14924 9660 15064
rect 3360 14896 3528 14924
rect 4032 14896 4340 14924
rect 5068 14896 5180 14924
rect 6300 14896 6356 14924
rect 6692 14896 6776 14924
rect 7728 14896 7840 14924
rect 8456 14896 8512 14924
rect 9212 14896 9380 14924
rect 3416 14868 3556 14896
rect 3948 14868 4284 14896
rect 5040 14868 5124 14896
rect 6300 14868 6384 14896
rect 6720 14868 6804 14896
rect 7644 14868 7784 14896
rect 8484 14868 8540 14896
rect 9184 14868 9352 14896
rect 3444 14840 3612 14868
rect 3892 14840 4228 14868
rect 4984 14840 5096 14868
rect 6328 14840 6384 14868
rect 6776 14840 6832 14868
rect 7560 14840 7700 14868
rect 8512 14840 8540 14868
rect 9072 14840 9324 14868
rect 3472 14812 3640 14840
rect 3808 14812 4172 14840
rect 4928 14812 5040 14840
rect 6356 14812 6412 14840
rect 6804 14812 6888 14840
rect 7504 14812 7616 14840
rect 3500 14784 3668 14812
rect 3752 14784 4116 14812
rect 4872 14784 4984 14812
rect 6356 14784 6440 14812
rect 6860 14784 6916 14812
rect 7420 14784 7532 14812
rect 3556 14756 4032 14784
rect 4816 14756 4928 14784
rect 6384 14756 6468 14784
rect 6888 14756 6972 14784
rect 7336 14756 7476 14784
rect 3584 14728 3976 14756
rect 4760 14728 4872 14756
rect 5404 14728 5460 14756
rect 6412 14728 6496 14756
rect 6916 14728 7000 14756
rect 7252 14728 7392 14756
rect 3612 14700 3920 14728
rect 4704 14700 4816 14728
rect 5432 14700 5488 14728
rect 6440 14700 6524 14728
rect 6972 14700 7056 14728
rect 7196 14700 7308 14728
rect 3640 14672 3864 14700
rect 4648 14672 4760 14700
rect 5320 14672 5404 14700
rect 5460 14672 5516 14700
rect 6468 14672 6552 14700
rect 7000 14672 7252 14700
rect 3696 14644 3836 14672
rect 4620 14644 4704 14672
rect 5264 14644 5348 14672
rect 5488 14644 5544 14672
rect 6524 14644 6580 14672
rect 3724 14616 3892 14644
rect 4564 14616 4648 14644
rect 5208 14616 5320 14644
rect 5516 14616 5572 14644
rect 6552 14616 6608 14644
rect 6944 14616 7028 14644
rect 3752 14588 3920 14616
rect 4508 14588 4592 14616
rect 5152 14588 5292 14616
rect 5544 14588 5600 14616
rect 6580 14588 6636 14616
rect 6860 14588 7140 14616
rect 3752 14560 3948 14588
rect 4452 14560 4536 14588
rect 4900 14560 4928 14588
rect 5124 14560 5320 14588
rect 5572 14560 5628 14588
rect 6804 14560 7196 14588
rect 3752 14532 3976 14560
rect 4396 14532 4480 14560
rect 4816 14532 4900 14560
rect 4928 14532 4956 14560
rect 5124 14532 5348 14560
rect 5600 14532 5656 14560
rect 6720 14532 7252 14560
rect 3752 14504 4004 14532
rect 4340 14504 4424 14532
rect 4760 14504 4844 14532
rect 4928 14504 4984 14532
rect 5152 14504 5376 14532
rect 5628 14504 5684 14532
rect 6664 14504 7308 14532
rect 3724 14476 4032 14504
rect 4284 14476 4368 14504
rect 4704 14476 4760 14504
rect 4956 14476 4984 14504
rect 5180 14476 5404 14504
rect 5656 14476 5712 14504
rect 6580 14476 7336 14504
rect 3724 14448 4088 14476
rect 4228 14448 4312 14476
rect 4648 14448 4704 14476
rect 4984 14448 5012 14476
rect 5180 14448 5432 14476
rect 5684 14448 5740 14476
rect 6524 14448 6748 14476
rect 6804 14448 7364 14476
rect 3696 14420 4116 14448
rect 4200 14420 4256 14448
rect 4592 14420 4648 14448
rect 5012 14420 5040 14448
rect 5208 14420 5460 14448
rect 5712 14420 5768 14448
rect 6468 14420 6692 14448
rect 6832 14420 7420 14448
rect 2632 14392 3248 14420
rect 3696 14392 4144 14420
rect 4592 14392 4620 14420
rect 5012 14392 5068 14420
rect 5236 14392 5460 14420
rect 5740 14392 5796 14420
rect 6384 14392 6636 14420
rect 6832 14392 7448 14420
rect 9044 14392 9072 14840
rect 9212 14812 9296 14840
rect 9240 14784 9268 14812
rect 9156 14700 9240 14728
rect 9156 14672 9184 14700
rect 9240 14672 9268 14700
rect 9632 14672 9660 14756
rect 9240 14644 9296 14672
rect 9268 14616 9296 14644
rect 9604 14616 9632 14672
rect 9296 14588 9324 14616
rect 9576 14588 9604 14616
rect 9324 14560 9352 14588
rect 9520 14560 9576 14588
rect 9352 14532 9408 14560
rect 9464 14532 9548 14560
rect 2464 14364 3388 14392
rect 3668 14364 4172 14392
rect 2380 14336 2660 14364
rect 3220 14336 3472 14364
rect 3668 14336 4004 14364
rect 4032 14336 4200 14364
rect 2268 14308 2520 14336
rect 3360 14308 3556 14336
rect 3640 14308 3976 14336
rect 4060 14308 4228 14336
rect 4564 14308 4592 14392
rect 4984 14364 5040 14392
rect 5264 14364 5488 14392
rect 5768 14364 5824 14392
rect 6328 14364 6552 14392
rect 6832 14364 7504 14392
rect 4928 14336 4984 14364
rect 5292 14336 5516 14364
rect 5796 14336 5852 14364
rect 6272 14336 6496 14364
rect 6720 14336 7532 14364
rect 4872 14308 4928 14336
rect 5320 14308 5544 14336
rect 5824 14308 5880 14336
rect 6272 14308 6440 14336
rect 6636 14308 6832 14336
rect 6888 14308 7560 14336
rect 2212 14280 2408 14308
rect 3444 14280 3976 14308
rect 4088 14280 4256 14308
rect 4564 14280 4620 14308
rect 4816 14280 4872 14308
rect 5348 14280 5572 14308
rect 5852 14280 5908 14308
rect 2128 14252 2324 14280
rect 3528 14252 3948 14280
rect 4144 14252 4284 14280
rect 4592 14252 4620 14280
rect 4732 14252 4816 14280
rect 5376 14252 5600 14280
rect 5880 14252 5936 14280
rect 6244 14252 6356 14308
rect 6552 14280 6664 14308
rect 6692 14280 6748 14308
rect 6888 14280 7616 14308
rect 6468 14252 6608 14280
rect 6776 14252 6832 14280
rect 6888 14252 7644 14280
rect 2072 14224 2240 14252
rect 3584 14224 3948 14252
rect 4172 14224 4312 14252
rect 4592 14224 4648 14252
rect 4676 14224 4760 14252
rect 5404 14224 5628 14252
rect 5908 14224 5964 14252
rect 6244 14224 6328 14252
rect 6412 14224 6552 14252
rect 6720 14224 6776 14252
rect 6888 14224 7532 14252
rect 7616 14224 7700 14252
rect 9072 14224 9100 14364
rect 9156 14280 9184 14532
rect 9828 14364 10024 14392
rect 9800 14336 9828 14364
rect 9996 14336 10052 14364
rect 10892 14336 11172 14364
rect 9772 14280 9800 14336
rect 10024 14308 10080 14336
rect 1988 14196 2156 14224
rect 1932 14168 2100 14196
rect 2492 14168 3136 14196
rect 3584 14168 3920 14224
rect 4200 14196 4340 14224
rect 4620 14196 4676 14224
rect 5404 14196 5656 14224
rect 5936 14196 5992 14224
rect 6244 14196 6468 14224
rect 6636 14196 6720 14224
rect 6832 14196 7476 14224
rect 7644 14196 7728 14224
rect 4228 14168 4368 14196
rect 5432 14168 5656 14196
rect 5964 14168 6020 14196
rect 1876 14140 2016 14168
rect 2380 14140 3276 14168
rect 3556 14140 3892 14168
rect 4256 14140 4396 14168
rect 5460 14140 5684 14168
rect 5992 14140 6020 14168
rect 6244 14168 6412 14196
rect 6552 14168 6664 14196
rect 6776 14168 6832 14196
rect 6944 14168 7392 14196
rect 7700 14168 7784 14196
rect 1820 14112 1960 14140
rect 2268 14112 2632 14140
rect 3108 14112 3360 14140
rect 3556 14112 3920 14140
rect 4284 14112 4424 14140
rect 5488 14112 5712 14140
rect 6020 14112 6048 14140
rect 6244 14112 6356 14168
rect 6468 14140 6608 14168
rect 6832 14140 6916 14168
rect 6944 14140 7336 14168
rect 7756 14140 7812 14168
rect 6384 14112 6552 14140
rect 6748 14112 6832 14140
rect 6944 14112 7280 14140
rect 7812 14112 7868 14140
rect 8596 14112 8652 14140
rect 9100 14112 9128 14224
rect 9184 14112 9212 14280
rect 9744 14252 9800 14280
rect 10052 14252 10080 14308
rect 10892 14308 11200 14336
rect 11452 14308 11592 14364
rect 10892 14280 11228 14308
rect 10892 14252 10976 14280
rect 11116 14252 11228 14280
rect 11424 14280 11592 14308
rect 11424 14252 11480 14280
rect 9604 14224 9772 14252
rect 9576 14196 9604 14224
rect 9548 14168 9604 14196
rect 9548 14140 9576 14168
rect 9660 14140 9800 14168
rect 1764 14084 1904 14112
rect 2184 14084 2492 14112
rect 3248 14084 3360 14112
rect 1736 14056 1848 14084
rect 2128 14056 2380 14084
rect 3332 14056 3360 14084
rect 3528 14084 3976 14112
rect 4312 14084 4452 14112
rect 5516 14084 5740 14112
rect 6048 14084 6076 14112
rect 6272 14084 6468 14112
rect 6664 14084 6776 14112
rect 6888 14084 6972 14112
rect 7000 14084 7196 14112
rect 7840 14084 7896 14112
rect 8512 14084 8596 14112
rect 8624 14084 8680 14112
rect 3528 14056 3864 14084
rect 3892 14056 4004 14084
rect 4340 14056 4480 14084
rect 5544 14056 5768 14084
rect 6048 14056 6104 14084
rect 6272 14056 6412 14084
rect 6608 14056 6720 14084
rect 6832 14056 6888 14084
rect 6972 14056 7000 14084
rect 7028 14056 7140 14084
rect 8456 14056 8540 14084
rect 1680 14028 1792 14056
rect 2044 14028 2296 14056
rect 1624 14000 1764 14028
rect 1988 14000 2212 14028
rect 3500 14000 3836 14056
rect 3948 14028 4060 14056
rect 4368 14028 4508 14056
rect 5572 14028 5796 14056
rect 6076 14028 6132 14056
rect 6272 14028 6384 14056
rect 6524 14028 6664 14056
rect 6888 14028 6972 14056
rect 7028 14028 7084 14056
rect 8400 14028 8540 14056
rect 8652 14028 8680 14084
rect 3976 14000 4088 14028
rect 4396 14000 4536 14028
rect 5600 14000 5824 14028
rect 6104 14000 6160 14028
rect 6300 14000 6412 14028
rect 6440 14000 6580 14028
rect 6804 14000 6888 14028
rect 1596 13972 1708 14000
rect 1960 13972 2156 14000
rect 1596 13944 1736 13972
rect 1904 13944 2100 13972
rect 3472 13944 3808 14000
rect 4004 13972 4116 14000
rect 4424 13972 4564 14000
rect 5600 13972 5852 14000
rect 6132 13972 6188 14000
rect 6300 13972 6524 14000
rect 6720 13972 6832 14000
rect 7056 13972 7084 14028
rect 8344 14000 8540 14028
rect 8316 13972 8568 14000
rect 8680 13972 8708 14028
rect 9128 14000 9156 14112
rect 4060 13944 4144 13972
rect 4452 13944 4592 13972
rect 5628 13944 5880 13972
rect 6160 13944 6216 13972
rect 6328 13944 6468 13972
rect 6664 13944 6776 13972
rect 6916 13944 6944 13972
rect 8260 13944 8316 13972
rect 1652 13916 2044 13944
rect 1708 13888 2016 13916
rect 3444 13888 3780 13944
rect 4088 13916 4172 13944
rect 4480 13916 4620 13944
rect 5656 13916 5880 13944
rect 6188 13916 6244 13944
rect 6356 13916 6468 13944
rect 6580 13916 6720 13944
rect 6888 13916 7112 13944
rect 8232 13916 8288 13944
rect 8372 13916 8568 13972
rect 8708 13916 8736 13972
rect 9156 13944 9184 14000
rect 9212 13972 9240 14112
rect 9520 14084 9548 14140
rect 9632 14112 9660 14140
rect 9772 14112 9828 14140
rect 9604 14084 9660 14112
rect 9800 14084 9828 14112
rect 9492 14056 9520 14084
rect 9604 14056 9632 14084
rect 9464 14000 9492 14056
rect 9576 14028 9604 14056
rect 9828 14028 9856 14084
rect 9548 14000 9604 14028
rect 9856 14000 9884 14028
rect 9436 13972 9464 14000
rect 9548 13972 9576 14000
rect 9856 13972 9912 14000
rect 9128 13916 9212 13944
rect 4116 13888 4200 13916
rect 4508 13888 4648 13916
rect 5684 13888 5908 13916
rect 6132 13888 6188 13916
rect 6216 13888 6272 13916
rect 6356 13888 6664 13916
rect 6972 13888 7140 13916
rect 8204 13888 8232 13916
rect 8372 13888 8596 13916
rect 1764 13860 2240 13888
rect 1708 13832 2520 13860
rect 3416 13832 3752 13888
rect 4144 13860 4228 13888
rect 4536 13860 4676 13888
rect 5712 13860 5936 13888
rect 6076 13860 6132 13888
rect 6244 13860 6580 13888
rect 7084 13860 7140 13888
rect 8176 13860 8204 13888
rect 4172 13832 4256 13860
rect 4564 13832 4704 13860
rect 5740 13832 5964 13860
rect 6020 13832 6104 13860
rect 6412 13832 6552 13860
rect 6664 13832 6692 13860
rect 7084 13832 7168 13860
rect 1680 13804 2632 13832
rect 1652 13776 2240 13804
rect 2436 13776 2716 13804
rect 3388 13776 3724 13832
rect 3976 13804 4004 13832
rect 4200 13804 4284 13832
rect 4592 13804 4732 13832
rect 5768 13804 6048 13832
rect 6440 13804 6580 13832
rect 3976 13776 4060 13804
rect 4228 13776 4312 13804
rect 4592 13776 4760 13804
rect 5796 13776 5992 13804
rect 6468 13776 6608 13804
rect 6692 13776 6720 13832
rect 7112 13804 7168 13832
rect 8148 13832 8204 13860
rect 8400 13860 8596 13888
rect 8736 13888 8764 13916
rect 8960 13888 9128 13916
rect 9156 13888 9212 13916
rect 9240 13888 9268 13972
rect 9408 13944 9464 13972
rect 9408 13916 9436 13944
rect 9520 13916 9548 13972
rect 9884 13944 9940 13972
rect 10080 13944 10108 14252
rect 10864 14224 10976 14252
rect 10864 14112 10948 14224
rect 11144 14196 11228 14252
rect 10836 13972 10920 14112
rect 11116 14056 11200 14196
rect 11396 14168 11480 14252
rect 11368 14084 11452 14168
rect 9912 13916 9968 13944
rect 10052 13916 10080 13944
rect 9380 13888 9408 13916
rect 9492 13888 9520 13916
rect 9968 13888 10052 13916
rect 8736 13860 8932 13888
rect 9184 13860 9268 13888
rect 8148 13804 8176 13832
rect 8400 13804 8624 13860
rect 9212 13832 9268 13860
rect 9352 13860 9408 13888
rect 9464 13860 9520 13888
rect 9576 13860 9632 13888
rect 10808 13860 10892 13972
rect 11088 13944 11172 14056
rect 11340 14028 11424 14084
rect 11508 14028 11592 14280
rect 11788 14252 11928 14364
rect 12096 14280 12180 14364
rect 11760 14196 11928 14252
rect 11760 14112 11844 14196
rect 11340 14000 11396 14028
rect 11508 14000 11564 14028
rect 11312 13944 11396 14000
rect 9352 13832 9632 13860
rect 9660 13832 9688 13860
rect 10780 13832 10892 13860
rect 11060 13916 11172 13944
rect 9240 13804 9296 13832
rect 9324 13804 9352 13832
rect 9520 13804 9576 13832
rect 9688 13804 9716 13832
rect 1624 13748 2184 13776
rect 2352 13748 2772 13776
rect 1596 13720 2128 13748
rect 2296 13720 2800 13748
rect 3360 13720 3696 13776
rect 4004 13748 4088 13776
rect 4256 13748 4340 13776
rect 4620 13748 4788 13776
rect 5824 13748 5936 13776
rect 6496 13748 6608 13776
rect 4032 13720 4116 13748
rect 4284 13720 4368 13748
rect 4648 13720 4816 13748
rect 1568 13692 2072 13720
rect 2240 13692 2856 13720
rect 1540 13664 2044 13692
rect 2184 13664 2632 13692
rect 2772 13664 2884 13692
rect 3332 13664 3668 13720
rect 4060 13692 4144 13720
rect 4312 13692 4396 13720
rect 4676 13692 4816 13720
rect 6524 13692 6636 13748
rect 6720 13720 6748 13776
rect 7112 13748 7196 13804
rect 7140 13720 7196 13748
rect 8120 13720 8148 13804
rect 8428 13748 8652 13804
rect 9240 13776 9324 13804
rect 9492 13776 9520 13804
rect 9716 13776 9744 13804
rect 9268 13748 9324 13776
rect 4088 13664 4172 13692
rect 4340 13664 4424 13692
rect 4704 13664 4844 13692
rect 6496 13664 6664 13692
rect 6748 13664 6776 13720
rect 7140 13692 7224 13720
rect 8456 13692 8680 13748
rect 9464 13720 9492 13776
rect 9660 13748 10136 13776
rect 9632 13720 9996 13748
rect 10136 13720 10164 13748
rect 10780 13720 10864 13832
rect 11060 13804 11144 13916
rect 11284 13860 11368 13944
rect 11032 13776 11144 13804
rect 11256 13832 11340 13860
rect 11480 13832 11564 14000
rect 11732 13972 11816 14112
rect 11704 13860 11788 13972
rect 11256 13776 11564 13832
rect 1512 13636 1988 13664
rect 2128 13636 2520 13664
rect 2828 13636 2912 13664
rect 1484 13608 1960 13636
rect 2072 13608 2436 13636
rect 2856 13608 2912 13636
rect 3304 13608 3640 13664
rect 4116 13636 4200 13664
rect 4368 13636 4452 13664
rect 4732 13636 4872 13664
rect 6440 13636 6496 13664
rect 6580 13636 6664 13664
rect 4144 13608 4228 13636
rect 4396 13608 4452 13636
rect 4760 13608 4900 13636
rect 6356 13608 6440 13636
rect 6580 13608 6692 13636
rect 1456 13580 1932 13608
rect 2044 13580 2352 13608
rect 2856 13580 2940 13608
rect 3304 13580 3612 13608
rect 4172 13580 4256 13608
rect 4396 13580 4480 13608
rect 4788 13580 4928 13608
rect 6300 13580 6384 13608
rect 6608 13580 6692 13608
rect 6776 13608 6804 13664
rect 7168 13636 7224 13692
rect 7168 13608 7252 13636
rect 8120 13608 8148 13692
rect 8484 13636 8708 13692
rect 8512 13608 8736 13636
rect 8792 13608 8820 13636
rect 9436 13608 9464 13720
rect 9604 13692 9996 13720
rect 6776 13580 6832 13608
rect 1456 13552 1876 13580
rect 2016 13552 2296 13580
rect 2884 13552 2968 13580
rect 1428 13524 1848 13552
rect 1960 13524 2240 13552
rect 2912 13524 2968 13552
rect 3276 13552 3612 13580
rect 4200 13552 4256 13580
rect 4424 13552 4508 13580
rect 4816 13552 4956 13580
rect 6244 13552 6328 13580
rect 3276 13524 3584 13552
rect 4200 13524 4284 13552
rect 4452 13524 4536 13552
rect 1400 13496 1820 13524
rect 1932 13496 2212 13524
rect 2912 13496 2996 13524
rect 1372 13468 1792 13496
rect 1904 13468 2156 13496
rect 1372 13440 1764 13468
rect 1876 13440 2128 13468
rect 1344 13412 1736 13440
rect 1848 13412 2072 13440
rect 2940 13412 2996 13496
rect 3248 13468 3584 13524
rect 4228 13496 4312 13524
rect 4480 13496 4536 13524
rect 4844 13524 4984 13552
rect 6160 13524 6272 13552
rect 6636 13524 6720 13580
rect 6804 13552 6832 13580
rect 7196 13552 7252 13608
rect 8148 13552 8176 13608
rect 8512 13580 8764 13608
rect 8540 13552 8708 13580
rect 9464 13552 9492 13608
rect 9576 13580 9968 13692
rect 10164 13580 10192 13720
rect 10752 13608 10836 13720
rect 11032 13664 11116 13776
rect 11228 13748 11564 13776
rect 11228 13692 11312 13748
rect 11004 13636 11088 13664
rect 11200 13636 11284 13692
rect 10976 13608 11088 13636
rect 11172 13608 11284 13636
rect 11480 13608 11564 13748
rect 11676 13832 11788 13860
rect 11676 13720 11760 13832
rect 10752 13580 11060 13608
rect 9604 13552 9996 13580
rect 10136 13552 10164 13580
rect 6804 13524 6860 13552
rect 4844 13496 5012 13524
rect 6104 13496 6216 13524
rect 6664 13496 6748 13524
rect 4256 13468 4340 13496
rect 4480 13468 4564 13496
rect 4872 13468 5040 13496
rect 6020 13468 6160 13496
rect 6636 13468 6748 13496
rect 6832 13468 6860 13524
rect 7224 13468 7280 13552
rect 8176 13524 8204 13552
rect 8540 13524 8652 13552
rect 9464 13524 9520 13552
rect 9632 13524 10024 13552
rect 10108 13524 10164 13552
rect 10724 13552 11032 13580
rect 11172 13552 11256 13608
rect 11452 13552 11564 13608
rect 11648 13580 11732 13720
rect 11872 13692 11928 14196
rect 12068 14252 12180 14280
rect 12320 14252 12404 14364
rect 12544 14336 12824 14364
rect 12544 14280 12796 14336
rect 12544 14252 12628 14280
rect 12908 14252 12992 14364
rect 13384 14280 13692 14364
rect 13804 14336 14084 14364
rect 13804 14280 14056 14336
rect 14140 14280 14448 14364
rect 13580 14252 13664 14280
rect 13804 14252 13888 14280
rect 14336 14252 14420 14280
rect 14532 14252 14672 14364
rect 14840 14280 14924 14364
rect 12068 14140 12152 14252
rect 12040 14112 12152 14140
rect 12292 14224 12404 14252
rect 12516 14224 12628 14252
rect 12880 14224 12992 14252
rect 12292 14112 12376 14224
rect 12516 14112 12600 14224
rect 12880 14112 12964 14224
rect 13552 14196 13636 14252
rect 13776 14224 13888 14252
rect 13524 14140 13608 14196
rect 12040 14000 12124 14112
rect 12012 13888 12096 14000
rect 12264 13972 12348 14112
rect 12488 14000 12572 14112
rect 12488 13972 12712 14000
rect 12852 13972 12936 14112
rect 13496 14084 13580 14140
rect 13776 14112 13860 14224
rect 14308 14196 14392 14252
rect 14504 14196 14672 14252
rect 14280 14140 14364 14196
rect 13468 14028 13552 14084
rect 13440 13972 13524 14028
rect 13748 14000 13832 14112
rect 14252 14084 14336 14140
rect 14504 14112 14588 14196
rect 14224 14028 14308 14084
rect 13748 13972 13972 14000
rect 14196 13972 14280 14028
rect 14476 13972 14560 14112
rect 11984 13860 12096 13888
rect 12236 13860 12320 13972
rect 12460 13916 12712 13972
rect 12460 13860 12544 13916
rect 12824 13860 12908 13972
rect 13412 13916 13496 13972
rect 13720 13916 13972 13972
rect 14168 13916 14252 13972
rect 13384 13860 13468 13916
rect 13720 13860 13804 13916
rect 14140 13860 14224 13916
rect 14448 13860 14532 13972
rect 11984 13720 12068 13860
rect 12208 13832 12320 13860
rect 12432 13832 12544 13860
rect 12796 13832 12908 13860
rect 12208 13720 12292 13832
rect 12432 13720 12516 13832
rect 12796 13720 12880 13832
rect 13356 13804 13440 13860
rect 13692 13832 13804 13860
rect 13328 13748 13412 13804
rect 13300 13720 13384 13748
rect 13692 13720 13776 13832
rect 14112 13804 14196 13860
rect 14420 13832 14532 13860
rect 14084 13748 14168 13804
rect 14056 13720 14140 13748
rect 14420 13720 14504 13832
rect 11956 13692 12040 13720
rect 11872 13608 12040 13692
rect 10724 13524 11004 13552
rect 11144 13524 11228 13552
rect 11452 13524 11536 13552
rect 11620 13524 11704 13580
rect 11872 13524 12012 13608
rect 12180 13580 12264 13720
rect 12404 13608 12488 13720
rect 12768 13608 12852 13720
rect 13272 13692 13384 13720
rect 13272 13664 13356 13692
rect 13244 13636 13356 13664
rect 13244 13608 13328 13636
rect 13664 13608 13748 13720
rect 14028 13692 14140 13720
rect 14028 13664 14112 13692
rect 14000 13636 14112 13664
rect 14000 13608 14084 13636
rect 12404 13580 12656 13608
rect 12768 13580 13020 13608
rect 12152 13524 12236 13580
rect 12376 13524 12656 13580
rect 12740 13524 12992 13580
rect 13216 13524 13524 13608
rect 13664 13580 13916 13608
rect 13636 13524 13916 13580
rect 13972 13524 14280 13608
rect 14392 13580 14476 13720
rect 14616 13692 14672 14196
rect 14812 14252 14924 14280
rect 15064 14252 15148 14364
rect 15372 14336 15568 14364
rect 15344 14308 15596 14336
rect 15288 14280 15596 14308
rect 15288 14252 15400 14280
rect 14812 14140 14896 14252
rect 14784 14112 14896 14140
rect 15036 14224 15148 14252
rect 15260 14224 15372 14252
rect 15036 14112 15120 14224
rect 15260 14140 15344 14224
rect 15232 14112 15344 14140
rect 15512 14196 15624 14280
rect 15736 14252 15820 14364
rect 16016 14336 16128 14364
rect 16016 14308 16100 14336
rect 15988 14280 16072 14308
rect 15708 14224 15820 14252
rect 15960 14252 16072 14280
rect 15960 14224 16044 14252
rect 14784 14000 14868 14112
rect 14756 13888 14840 14000
rect 15008 13972 15092 14112
rect 15232 14000 15316 14112
rect 15512 14084 15596 14196
rect 15708 14112 15792 14224
rect 15932 14168 16016 14224
rect 15904 14140 15988 14168
rect 15876 14112 15988 14140
rect 15484 14056 15568 14084
rect 15680 14000 15764 14112
rect 15876 14084 15960 14112
rect 15848 14028 15932 14084
rect 15820 14000 15904 14028
rect 14728 13860 14840 13888
rect 14980 13860 15064 13972
rect 15204 13860 15288 14000
rect 15680 13972 15876 14000
rect 15652 13916 15876 13972
rect 15652 13860 15736 13916
rect 14728 13720 14812 13860
rect 14952 13832 15064 13860
rect 14952 13720 15036 13832
rect 15176 13748 15260 13860
rect 15624 13832 15736 13860
rect 15792 13860 15876 13916
rect 15148 13720 15260 13748
rect 15428 13804 15540 13832
rect 14700 13692 14784 13720
rect 14616 13608 14784 13692
rect 14364 13524 14448 13580
rect 14616 13524 14756 13608
rect 14924 13580 15008 13720
rect 15148 13636 15232 13720
rect 15428 13692 15512 13804
rect 15624 13720 15708 13832
rect 15792 13804 15904 13860
rect 15820 13720 15904 13804
rect 15400 13664 15512 13692
rect 15400 13636 15484 13664
rect 15148 13608 15260 13636
rect 15372 13608 15484 13636
rect 15148 13580 15456 13608
rect 15596 13580 15680 13720
rect 15820 13664 15932 13720
rect 15848 13580 15932 13664
rect 14896 13524 14980 13580
rect 15176 13552 15428 13580
rect 15204 13524 15400 13552
rect 15568 13524 15652 13580
rect 15848 13524 15960 13580
rect 8176 13496 8232 13524
rect 8512 13496 8596 13524
rect 9492 13496 9548 13524
rect 9660 13496 9716 13524
rect 9996 13496 10024 13524
rect 8204 13468 8260 13496
rect 8428 13468 8512 13496
rect 9548 13468 9660 13496
rect 3220 13412 3556 13468
rect 4284 13440 4368 13468
rect 4508 13440 4592 13468
rect 4900 13440 5040 13468
rect 5936 13440 6104 13468
rect 6608 13440 6636 13468
rect 4312 13412 4396 13440
rect 1316 13356 1708 13412
rect 1820 13384 2044 13412
rect 1792 13356 2016 13384
rect 2940 13356 3024 13412
rect 3192 13356 3528 13412
rect 4340 13384 4396 13412
rect 4536 13384 4620 13440
rect 4928 13412 5068 13440
rect 5852 13412 6048 13440
rect 6580 13412 6636 13440
rect 6692 13412 6776 13468
rect 6860 13412 6888 13468
rect 7252 13412 7308 13468
rect 8260 13440 8456 13468
rect 8848 13440 9128 13468
rect 9576 13440 9632 13468
rect 8316 13412 8400 13440
rect 8792 13412 8876 13440
rect 9072 13412 9576 13440
rect 4956 13384 5096 13412
rect 5768 13384 5964 13412
rect 6552 13384 6608 13412
rect 6720 13384 6804 13412
rect 4340 13356 4424 13384
rect 4564 13356 4648 13384
rect 4984 13356 5124 13384
rect 5684 13356 5908 13384
rect 6524 13356 6580 13384
rect 6748 13356 6804 13384
rect 6888 13356 6916 13412
rect 7280 13384 7308 13412
rect 8260 13384 8344 13412
rect 8736 13384 8820 13412
rect 9464 13384 9576 13412
rect 1288 13328 1680 13356
rect 1288 13300 1652 13328
rect 1764 13300 1988 13356
rect 2968 13328 3024 13356
rect 2716 13300 3024 13328
rect 3164 13300 3500 13356
rect 4368 13328 4452 13356
rect 4396 13300 4452 13328
rect 4592 13328 4648 13356
rect 5012 13328 5152 13356
rect 5600 13328 5852 13356
rect 6496 13328 6552 13356
rect 6748 13328 6832 13356
rect 6888 13328 6944 13356
rect 7280 13328 7336 13384
rect 8232 13356 8288 13384
rect 8708 13356 8764 13384
rect 9576 13356 9632 13384
rect 8064 13328 8232 13356
rect 8652 13328 8708 13356
rect 9604 13328 9660 13356
rect 4592 13300 4676 13328
rect 5012 13300 5180 13328
rect 5488 13300 5768 13328
rect 6496 13300 6524 13328
rect 1260 13272 1624 13300
rect 1736 13272 1960 13300
rect 2604 13272 2828 13300
rect 2884 13272 3024 13300
rect 1232 13244 1624 13272
rect 1708 13244 1960 13272
rect 2520 13244 2660 13272
rect 2968 13244 3024 13272
rect 3136 13272 3584 13300
rect 4396 13272 4480 13300
rect 4620 13272 4704 13300
rect 5040 13272 5180 13300
rect 5404 13272 5684 13300
rect 6468 13272 6524 13300
rect 6776 13300 6832 13328
rect 6916 13300 6944 13328
rect 6776 13272 6860 13300
rect 6916 13272 6972 13300
rect 7308 13272 7364 13328
rect 7868 13300 8092 13328
rect 8176 13300 8232 13328
rect 8596 13300 8652 13328
rect 9660 13300 9716 13328
rect 7812 13272 7952 13300
rect 8008 13272 8036 13300
rect 3136 13244 3668 13272
rect 4424 13244 4508 13272
rect 4648 13244 4704 13272
rect 5068 13244 5208 13272
rect 5292 13244 5628 13272
rect 6440 13244 6496 13272
rect 6804 13244 6860 13272
rect 6944 13244 6972 13272
rect 7336 13244 7364 13272
rect 7784 13244 7812 13272
rect 7840 13244 7952 13272
rect 1232 13188 1596 13244
rect 1680 13188 1960 13244
rect 2464 13216 2576 13244
rect 2940 13216 3024 13244
rect 2408 13188 2492 13216
rect 1204 13160 1568 13188
rect 1652 13160 1960 13188
rect 2352 13160 2436 13188
rect 1204 13132 1540 13160
rect 1652 13132 1988 13160
rect 2324 13132 2408 13160
rect 2940 13132 2996 13216
rect 3108 13188 3444 13244
rect 3528 13216 3752 13244
rect 3612 13188 3808 13216
rect 4452 13188 4536 13244
rect 4648 13216 4732 13244
rect 5096 13216 5544 13244
rect 6412 13216 6468 13244
rect 6804 13216 6888 13244
rect 6944 13216 7000 13244
rect 4676 13188 4732 13216
rect 5124 13188 5460 13216
rect 6384 13188 6440 13216
rect 6832 13188 6888 13216
rect 6972 13188 7000 13216
rect 7336 13188 7392 13244
rect 3080 13132 3416 13188
rect 3696 13160 3920 13188
rect 4480 13160 4564 13188
rect 4676 13160 4760 13188
rect 5124 13160 5376 13188
rect 6356 13160 6412 13188
rect 6832 13160 6916 13188
rect 6972 13160 7028 13188
rect 3780 13132 4004 13160
rect 4508 13132 4564 13160
rect 4704 13132 4760 13160
rect 5152 13132 5292 13160
rect 6328 13132 6384 13160
rect 6860 13132 6916 13160
rect 7000 13132 7028 13160
rect 7364 13160 7392 13188
rect 7756 13160 7784 13244
rect 7364 13132 7420 13160
rect 7840 13132 7924 13244
rect 1176 13104 1540 13132
rect 1624 13104 1988 13132
rect 2296 13104 2352 13132
rect 1176 13048 1512 13104
rect 1148 13020 1512 13048
rect 1596 13076 2016 13104
rect 2268 13076 2324 13104
rect 2912 13076 2996 13132
rect 3052 13104 3416 13132
rect 3556 13104 3584 13132
rect 3808 13104 4088 13132
rect 4508 13104 4592 13132
rect 4704 13104 4788 13132
rect 3052 13076 3584 13104
rect 3780 13076 4172 13104
rect 4536 13076 4620 13104
rect 1596 13048 2044 13076
rect 2240 13048 2296 13076
rect 1596 13020 2100 13048
rect 2212 13020 2268 13048
rect 2912 13020 3360 13076
rect 3416 13048 3612 13076
rect 3752 13048 4284 13076
rect 4564 13048 4620 13076
rect 4732 13076 4788 13104
rect 5152 13104 5236 13132
rect 6300 13104 6356 13132
rect 6860 13104 6944 13132
rect 7000 13104 7056 13132
rect 7392 13104 7420 13132
rect 3444 13020 3612 13048
rect 3724 13020 4368 13048
rect 4564 13020 4648 13048
rect 4732 13020 4816 13076
rect 5152 13048 5264 13104
rect 6272 13076 6328 13104
rect 6888 13076 6944 13104
rect 7028 13076 7056 13104
rect 6244 13048 6300 13076
rect 6888 13048 6972 13076
rect 1148 12964 1484 13020
rect 1568 12992 2240 13020
rect 1568 12964 2212 12992
rect 2996 12964 3332 13020
rect 3416 12992 3640 13020
rect 3696 12992 4144 13020
rect 4228 12992 4508 13020
rect 4592 12992 4816 13020
rect 5180 12992 5292 13048
rect 6216 13020 6272 13048
rect 6188 12992 6244 13020
rect 6916 12992 6972 13048
rect 7028 13020 7084 13076
rect 7056 12992 7084 13020
rect 3416 12964 3808 12992
rect 3892 12964 4172 12992
rect 1120 12880 1456 12964
rect 1540 12936 2184 12964
rect 2772 12936 2940 12964
rect 2968 12936 3304 12964
rect 1540 12908 1708 12936
rect 1820 12908 2184 12936
rect 2660 12908 3304 12936
rect 1540 12880 1680 12908
rect 1932 12880 2156 12908
rect 2604 12880 2828 12908
rect 2912 12880 3276 12908
rect 1092 12768 1428 12880
rect 1512 12824 1680 12880
rect 2044 12852 2128 12880
rect 2548 12852 2688 12880
rect 2716 12852 2828 12880
rect 2940 12852 3276 12880
rect 3388 12852 3780 12964
rect 3948 12936 4172 12964
rect 4004 12908 4172 12936
rect 4256 12964 4760 12992
rect 5208 12964 5320 12992
rect 6160 12964 6216 12992
rect 4256 12936 4704 12964
rect 5208 12936 5348 12964
rect 6104 12936 6188 12964
rect 6944 12936 7000 12992
rect 7056 12964 7112 12992
rect 7084 12936 7112 12964
rect 4256 12908 4592 12936
rect 5236 12908 5348 12936
rect 6076 12908 6160 12936
rect 2072 12824 2128 12852
rect 2520 12824 2632 12852
rect 1512 12796 1652 12824
rect 2072 12796 2100 12824
rect 2492 12796 2576 12824
rect 1092 12740 1400 12768
rect 1064 12600 1400 12740
rect 1484 12712 1652 12796
rect 2044 12768 2100 12796
rect 2464 12768 2548 12796
rect 2744 12768 2828 12852
rect 2912 12796 3248 12852
rect 2884 12768 3248 12796
rect 3388 12824 3752 12852
rect 4032 12824 4200 12908
rect 2044 12740 2072 12768
rect 2436 12740 2520 12768
rect 2744 12740 2856 12768
rect 2884 12740 3276 12768
rect 3388 12740 3780 12824
rect 4060 12740 4228 12824
rect 4284 12796 4620 12908
rect 1484 12656 1624 12712
rect 1064 12292 1372 12600
rect 1456 12404 1624 12656
rect 2016 12684 2072 12740
rect 2408 12712 2492 12740
rect 2408 12684 2464 12712
rect 2016 12628 2044 12684
rect 2380 12656 2464 12684
rect 2772 12684 3192 12740
rect 3220 12712 3304 12740
rect 3248 12684 3332 12712
rect 3388 12684 3808 12740
rect 4088 12684 4228 12740
rect 4312 12768 4620 12796
rect 2380 12628 2436 12656
rect 2772 12628 3164 12684
rect 3276 12656 3332 12684
rect 3416 12656 3864 12684
rect 3276 12628 3360 12656
rect 1988 12544 2044 12628
rect 2352 12600 2436 12628
rect 2352 12572 2408 12600
rect 2800 12572 3136 12628
rect 3304 12572 3360 12628
rect 3416 12572 3892 12656
rect 2352 12544 2492 12572
rect 1456 12376 1680 12404
rect 1456 12348 1764 12376
rect 1988 12348 2016 12544
rect 2324 12516 2688 12544
rect 2772 12516 3108 12572
rect 3304 12544 3388 12572
rect 2324 12488 3080 12516
rect 1456 12320 1876 12348
rect 1456 12292 1960 12320
rect 1988 12292 2044 12348
rect 2324 12320 2380 12488
rect 2436 12460 3080 12488
rect 2632 12432 3080 12460
rect 2744 12404 3248 12432
rect 3332 12404 3388 12544
rect 3444 12544 3892 12572
rect 4088 12544 4256 12684
rect 4312 12656 4648 12768
rect 3444 12488 3864 12544
rect 3472 12432 3864 12488
rect 2744 12348 3388 12404
rect 2744 12320 3024 12348
rect 3220 12320 3388 12348
rect 2324 12292 2408 12320
rect 2744 12292 2996 12320
rect 3332 12292 3388 12320
rect 3500 12292 3836 12432
rect 4116 12348 4256 12544
rect 1064 12180 1400 12292
rect 1456 12264 2044 12292
rect 1092 12124 1400 12180
rect 1484 12236 2044 12264
rect 2352 12236 2408 12292
rect 2716 12264 2996 12292
rect 2688 12236 2996 12264
rect 3304 12264 3388 12292
rect 3528 12264 3808 12292
rect 1484 12180 2072 12236
rect 2352 12208 2436 12236
rect 2660 12208 2800 12236
rect 1484 12152 1904 12180
rect 1988 12152 2072 12180
rect 2380 12180 2436 12208
rect 2632 12180 2772 12208
rect 2912 12180 3024 12236
rect 3304 12208 3360 12264
rect 3528 12236 3780 12264
rect 3584 12208 3752 12236
rect 4088 12208 4256 12348
rect 4340 12236 4648 12656
rect 5264 12628 5348 12908
rect 6048 12880 6132 12908
rect 6972 12880 7028 12936
rect 7084 12908 7140 12936
rect 6020 12852 6104 12880
rect 7000 12852 7028 12880
rect 7112 12880 7140 12908
rect 7112 12852 7168 12880
rect 5992 12824 6076 12852
rect 7000 12824 7056 12852
rect 7140 12824 7168 12852
rect 7728 12824 7756 13132
rect 7812 13020 7924 13132
rect 5964 12796 6048 12824
rect 7028 12796 7056 12824
rect 5936 12768 6020 12796
rect 5880 12740 5992 12768
rect 7028 12740 7084 12796
rect 5852 12712 5964 12740
rect 5824 12684 5936 12712
rect 5796 12656 5880 12684
rect 7056 12656 7084 12740
rect 5740 12628 5852 12656
rect 7056 12628 7112 12656
rect 5236 12572 5348 12628
rect 5712 12600 5824 12628
rect 7084 12600 7112 12628
rect 5684 12572 5796 12600
rect 7084 12572 7140 12600
rect 5236 12488 5320 12572
rect 5656 12544 5740 12572
rect 7112 12544 7168 12572
rect 5600 12516 5712 12544
rect 6524 12516 6552 12544
rect 7140 12516 7196 12544
rect 7728 12516 7756 12796
rect 7812 12544 7896 13020
rect 7980 12964 8008 13244
rect 8008 12880 8036 12964
rect 8064 12936 8092 13300
rect 8232 13272 8260 13300
rect 8540 13272 8596 13300
rect 8260 13244 8288 13272
rect 8512 13244 8540 13272
rect 9464 13244 9492 13300
rect 9716 13272 9772 13300
rect 10668 13272 15988 13328
rect 9716 13244 9828 13272
rect 10668 13244 15960 13272
rect 8260 13216 8316 13244
rect 9436 13216 9464 13244
rect 9716 13216 9856 13244
rect 8288 13188 8316 13216
rect 8596 13188 8652 13216
rect 9380 13188 9436 13216
rect 8316 13160 8344 13188
rect 8540 13160 8596 13188
rect 8652 13160 8708 13188
rect 9296 13160 9436 13188
rect 9716 13188 9912 13216
rect 10640 13188 15932 13244
rect 9716 13160 9940 13188
rect 8344 13048 8372 13160
rect 8540 13132 8568 13160
rect 8708 13132 8736 13160
rect 9296 13132 9324 13160
rect 8736 13104 8792 13132
rect 8540 13076 8568 13104
rect 8792 13076 8820 13104
rect 9324 13076 9352 13132
rect 9380 13104 9408 13160
rect 9716 13132 9996 13160
rect 10612 13132 15904 13188
rect 9688 13104 10024 13132
rect 10612 13104 15876 13132
rect 9408 13076 9464 13104
rect 9688 13076 10052 13104
rect 8540 13048 8596 13076
rect 8820 13048 8848 13076
rect 9296 13048 9352 13076
rect 9464 13048 9548 13076
rect 9660 13048 9716 13076
rect 9744 13048 10080 13076
rect 8316 12936 8372 13048
rect 8512 13020 8624 13048
rect 8484 12992 8652 13020
rect 8848 12992 8876 13048
rect 9212 13020 9296 13048
rect 9520 13020 9604 13048
rect 9660 13020 9688 13048
rect 9828 13020 10080 13048
rect 9156 12992 9240 13020
rect 9604 12992 9660 13020
rect 9884 12992 10080 13020
rect 8484 12964 8708 12992
rect 9100 12964 9156 12992
rect 9940 12964 10080 12992
rect 8456 12936 8764 12964
rect 8792 12936 8848 12964
rect 9044 12936 9100 12964
rect 9548 12936 9744 12964
rect 9996 12936 10052 12964
rect 8288 12908 8316 12936
rect 8260 12880 8288 12908
rect 8008 12852 8064 12880
rect 8036 12824 8064 12852
rect 8092 12824 8120 12880
rect 8232 12852 8288 12880
rect 8372 12880 8400 12936
rect 8456 12908 8792 12936
rect 8428 12880 8736 12908
rect 9044 12880 9072 12936
rect 9436 12908 9912 12936
rect 9352 12880 9996 12908
rect 8372 12852 8736 12880
rect 8204 12824 8260 12852
rect 8372 12824 8708 12852
rect 8064 12796 8204 12824
rect 8372 12796 8680 12824
rect 9016 12796 9044 12880
rect 9296 12852 9632 12880
rect 9716 12852 10080 12880
rect 9240 12824 9492 12852
rect 9884 12824 10164 12852
rect 9212 12796 9408 12824
rect 9968 12796 10220 12824
rect 8344 12768 8680 12796
rect 8736 12768 8764 12796
rect 8344 12740 8652 12768
rect 8316 12712 8652 12740
rect 8708 12740 8820 12768
rect 8988 12740 9016 12796
rect 9184 12768 9324 12796
rect 10052 12768 10276 12796
rect 9156 12740 9296 12768
rect 10136 12740 10332 12768
rect 8708 12712 8876 12740
rect 8960 12712 9016 12740
rect 9128 12712 9240 12740
rect 10192 12712 10388 12740
rect 8288 12684 8624 12712
rect 8680 12684 8904 12712
rect 8960 12684 8988 12712
rect 8288 12656 8596 12684
rect 8680 12656 8988 12684
rect 9100 12656 9212 12712
rect 9380 12684 9408 12712
rect 10248 12684 10444 12712
rect 9324 12656 9380 12684
rect 10304 12656 10472 12684
rect 8260 12628 8596 12656
rect 8652 12628 8960 12656
rect 8232 12600 8568 12628
rect 8624 12600 8960 12628
rect 9072 12628 9184 12656
rect 9296 12628 9352 12656
rect 10108 12628 10164 12656
rect 10360 12628 10528 12656
rect 9072 12600 9156 12628
rect 8232 12572 8540 12600
rect 8624 12572 8932 12600
rect 8204 12544 8540 12572
rect 8596 12544 8932 12572
rect 5572 12488 5684 12516
rect 5208 12404 5320 12488
rect 5544 12460 5628 12488
rect 6496 12460 6580 12516
rect 5488 12432 5600 12460
rect 5880 12432 5908 12460
rect 6468 12432 6552 12460
rect 7756 12432 7784 12516
rect 7812 12460 7924 12544
rect 8204 12516 8512 12544
rect 8176 12488 8512 12516
rect 8568 12516 8932 12544
rect 9044 12572 9156 12600
rect 9268 12600 9324 12628
rect 10136 12600 10192 12628
rect 10416 12600 10584 12628
rect 9268 12572 9296 12600
rect 10192 12572 10248 12600
rect 10472 12572 10612 12600
rect 8568 12488 8960 12516
rect 8148 12460 8484 12488
rect 8540 12460 9016 12488
rect 9044 12460 9128 12572
rect 5460 12404 5544 12432
rect 5852 12404 5908 12432
rect 5208 12376 5292 12404
rect 5432 12376 5516 12404
rect 5852 12376 5880 12404
rect 5964 12376 6048 12432
rect 6440 12404 6496 12432
rect 7784 12404 7812 12432
rect 7840 12404 7924 12460
rect 8120 12432 8456 12460
rect 8540 12432 9128 12460
rect 8092 12404 8456 12432
rect 8512 12404 9128 12432
rect 6440 12376 6468 12404
rect 6720 12376 6776 12404
rect 7784 12376 7924 12404
rect 8036 12376 8428 12404
rect 5180 12320 5292 12376
rect 5572 12348 5656 12376
rect 5824 12348 5880 12376
rect 5936 12348 6020 12376
rect 6664 12348 6804 12376
rect 7812 12348 8036 12376
rect 8092 12348 8400 12376
rect 8484 12348 9128 12404
rect 9240 12544 9296 12572
rect 10220 12544 10304 12572
rect 10500 12544 10668 12572
rect 9240 12376 9268 12544
rect 10276 12516 10332 12544
rect 10556 12516 10696 12544
rect 9800 12488 9940 12516
rect 10332 12488 10388 12516
rect 10612 12488 10752 12516
rect 9716 12460 9996 12488
rect 10360 12460 10416 12488
rect 10640 12460 10780 12488
rect 9688 12432 10052 12460
rect 10416 12432 10472 12460
rect 10696 12432 10808 12460
rect 9660 12404 9772 12432
rect 9968 12404 10080 12432
rect 10444 12404 10528 12432
rect 10724 12404 10864 12432
rect 9660 12376 9744 12404
rect 9828 12376 9912 12404
rect 9996 12376 10080 12404
rect 10500 12376 10556 12404
rect 10780 12376 10892 12404
rect 5572 12320 5684 12348
rect 5796 12320 5852 12348
rect 5936 12320 5964 12348
rect 6244 12320 6300 12348
rect 6608 12320 6804 12348
rect 7896 12320 7952 12348
rect 8064 12320 8400 12348
rect 8456 12320 9156 12348
rect 9240 12320 9296 12376
rect 9632 12348 9716 12376
rect 9772 12348 9968 12376
rect 9632 12320 9688 12348
rect 5180 12292 5264 12320
rect 5544 12292 5656 12320
rect 5152 12236 5264 12292
rect 5516 12264 5656 12292
rect 5768 12264 5824 12320
rect 6188 12292 6328 12320
rect 6384 12292 6468 12320
rect 6552 12292 6776 12320
rect 5880 12264 5936 12292
rect 6048 12264 6132 12292
rect 6160 12264 6300 12292
rect 6356 12264 6468 12292
rect 6524 12264 6664 12292
rect 6692 12264 6748 12292
rect 8036 12264 8372 12320
rect 8428 12264 9156 12320
rect 9268 12292 9296 12320
rect 9268 12264 9324 12292
rect 5488 12236 5656 12264
rect 5740 12236 5796 12264
rect 5852 12236 5936 12264
rect 6020 12236 6300 12264
rect 6328 12236 6440 12264
rect 6496 12236 6608 12264
rect 6664 12236 6748 12264
rect 8008 12236 8344 12264
rect 3276 12180 3360 12208
rect 2380 12152 2464 12180
rect 2604 12152 2744 12180
rect 2940 12152 3024 12180
rect 3248 12152 3332 12180
rect 3640 12152 3696 12208
rect 4088 12180 4228 12208
rect 1484 12124 1820 12152
rect 1092 12040 1428 12124
rect 1484 12096 1792 12124
rect 2044 12096 2100 12152
rect 2408 12096 2492 12152
rect 2576 12124 2716 12152
rect 2940 12124 3052 12152
rect 3248 12124 3304 12152
rect 3640 12124 3668 12152
rect 2548 12096 2688 12124
rect 2968 12096 3052 12124
rect 3220 12096 3304 12124
rect 3612 12096 3668 12124
rect 4060 12096 4228 12180
rect 4312 12124 4648 12236
rect 5124 12180 5236 12236
rect 5460 12208 5656 12236
rect 5712 12208 5936 12236
rect 5992 12208 6272 12236
rect 5460 12180 5516 12208
rect 5124 12152 5208 12180
rect 5432 12152 5488 12180
rect 5544 12152 5628 12208
rect 5712 12180 5908 12208
rect 5936 12180 6272 12208
rect 6300 12208 6580 12236
rect 6608 12208 6748 12236
rect 6832 12208 6916 12236
rect 6300 12180 6524 12208
rect 6580 12180 6720 12208
rect 6804 12180 6916 12208
rect 7980 12180 8316 12236
rect 8400 12208 9184 12264
rect 9296 12236 9324 12264
rect 9296 12208 9352 12236
rect 8372 12180 9184 12208
rect 9324 12180 9352 12208
rect 9604 12180 9688 12320
rect 9744 12264 9996 12348
rect 10024 12320 10108 12376
rect 10528 12348 10612 12376
rect 10808 12348 10948 12376
rect 10584 12320 10640 12348
rect 10836 12320 10976 12348
rect 9716 12236 9996 12264
rect 9744 12180 9996 12236
rect 10052 12208 10136 12320
rect 10640 12292 10696 12320
rect 10892 12292 11004 12320
rect 10668 12264 10752 12292
rect 10920 12264 11032 12292
rect 10724 12236 10780 12264
rect 10976 12236 11088 12264
rect 10752 12208 10836 12236
rect 11004 12208 11116 12236
rect 10052 12180 10108 12208
rect 10808 12180 10864 12208
rect 11032 12180 11144 12208
rect 5684 12152 5768 12180
rect 5796 12152 5964 12180
rect 5992 12152 6104 12180
rect 6132 12152 6244 12180
rect 6272 12152 6496 12180
rect 6552 12152 6860 12180
rect 7952 12152 8288 12180
rect 5096 12124 5208 12152
rect 5404 12124 5488 12152
rect 4312 12096 4620 12124
rect 1120 12012 1428 12040
rect 1512 12068 1792 12096
rect 2072 12068 2100 12096
rect 2436 12068 2660 12096
rect 2968 12068 3080 12096
rect 3192 12068 3276 12096
rect 3612 12068 3640 12096
rect 4060 12068 4200 12096
rect 1512 12012 1764 12068
rect 2072 12040 2128 12068
rect 2464 12040 2632 12068
rect 2996 12040 3080 12068
rect 3164 12040 3248 12068
rect 3584 12040 3640 12068
rect 1120 11928 1456 12012
rect 1540 11928 1736 12012
rect 2100 11984 2156 12040
rect 2492 12012 2604 12040
rect 2996 12012 3220 12040
rect 3584 12012 3612 12040
rect 2520 11984 2632 12012
rect 3024 11984 3192 12012
rect 3556 11984 3612 12012
rect 4032 11984 4200 12068
rect 4284 12012 4620 12096
rect 5068 12068 5180 12124
rect 5376 12096 5488 12124
rect 5516 12124 5628 12152
rect 5376 12068 5460 12096
rect 5040 12012 5152 12068
rect 5348 12012 5460 12068
rect 5516 12040 5600 12124
rect 5656 12096 5740 12152
rect 5796 12124 5936 12152
rect 5964 12124 6076 12152
rect 6104 12124 6216 12152
rect 6272 12124 6776 12152
rect 5768 12096 5908 12124
rect 5936 12096 6048 12124
rect 6104 12096 6356 12124
rect 5628 12068 5712 12096
rect 5740 12068 5880 12096
rect 5936 12068 6020 12096
rect 6076 12068 6356 12096
rect 6384 12096 6552 12124
rect 6608 12096 6720 12124
rect 7924 12096 8260 12152
rect 8344 12124 9212 12180
rect 9324 12124 9380 12180
rect 9632 12124 9716 12180
rect 9772 12152 9968 12180
rect 9800 12124 9940 12152
rect 10024 12124 10108 12180
rect 10836 12152 10920 12180
rect 11060 12152 11172 12180
rect 10892 12124 10948 12152
rect 11116 12124 11228 12152
rect 8316 12096 9240 12124
rect 9352 12096 9408 12124
rect 6384 12068 6524 12096
rect 6608 12068 6664 12096
rect 5628 12040 5852 12068
rect 5908 12040 6020 12068
rect 6104 12040 6188 12068
rect 6216 12040 6328 12068
rect 7896 12040 8232 12096
rect 8288 12068 9240 12096
rect 9380 12068 9408 12096
rect 9660 12096 9744 12124
rect 9996 12096 10080 12124
rect 10920 12096 11004 12124
rect 11144 12096 11256 12124
rect 9660 12068 9800 12096
rect 9940 12068 10052 12096
rect 10948 12068 11032 12096
rect 11172 12068 11284 12096
rect 8288 12040 9268 12068
rect 9380 12040 9436 12068
rect 9688 12040 10024 12068
rect 11004 12040 11088 12068
rect 11200 12040 11312 12068
rect 5488 12012 5684 12040
rect 5712 12012 5824 12040
rect 5936 12012 5992 12040
rect 6188 12012 6300 12040
rect 7868 12012 8204 12040
rect 8260 12012 9268 12040
rect 9408 12012 9436 12040
rect 9744 12012 9996 12040
rect 11032 12012 11116 12040
rect 11256 12012 11340 12040
rect 2128 11956 2184 11984
rect 2576 11956 2716 11984
rect 2996 11956 3164 11984
rect 1148 11872 1484 11928
rect 1568 11872 1736 11928
rect 2156 11900 2212 11956
rect 2604 11928 3108 11956
rect 3528 11928 3584 11984
rect 4004 11928 4172 11984
rect 4256 11928 4592 12012
rect 5012 11984 5124 12012
rect 4984 11956 5096 11984
rect 2688 11900 3052 11928
rect 3500 11900 3556 11928
rect 2184 11872 2240 11900
rect 3472 11872 3556 11900
rect 3976 11872 4144 11928
rect 1148 11844 1512 11872
rect 1176 11816 1512 11844
rect 1596 11844 1764 11872
rect 2212 11844 2268 11872
rect 3444 11844 3584 11872
rect 1596 11816 1792 11844
rect 2240 11816 2296 11844
rect 3416 11816 3584 11844
rect 3948 11844 4144 11872
rect 4228 11900 4592 11928
rect 4956 11928 5096 11956
rect 5320 11956 5432 12012
rect 5488 11956 5656 12012
rect 5740 11984 5768 12012
rect 6160 11984 6300 12012
rect 6132 11956 6272 11984
rect 6776 11956 6804 11984
rect 7840 11956 8176 12012
rect 8260 11984 9296 12012
rect 9408 11984 9464 12012
rect 9828 11984 9912 12012
rect 11088 11984 11144 12012
rect 11284 11984 11368 12012
rect 8232 11956 9324 11984
rect 5320 11928 5404 11956
rect 5488 11928 5628 11956
rect 6104 11928 6216 11956
rect 6720 11928 6748 11956
rect 7812 11928 8148 11956
rect 8204 11928 9324 11956
rect 9436 11956 9464 11984
rect 11116 11956 11200 11984
rect 11312 11956 11424 11984
rect 9436 11928 9492 11956
rect 11144 11928 11228 11956
rect 11340 11928 11452 11956
rect 12964 11928 13048 11956
rect 4956 11900 5124 11928
rect 5320 11900 5376 11928
rect 5488 11900 5600 11928
rect 6076 11900 6132 11928
rect 6664 11900 6692 11928
rect 4228 11844 4564 11900
rect 4956 11872 5208 11900
rect 6048 11872 6104 11900
rect 6580 11872 6636 11900
rect 7784 11872 8120 11928
rect 8204 11900 9352 11928
rect 9464 11900 9492 11928
rect 11200 11900 11284 11928
rect 11368 11900 11480 11928
rect 8176 11872 8960 11900
rect 9156 11872 9380 11900
rect 9464 11872 9520 11900
rect 11228 11872 11312 11900
rect 11424 11872 11508 11900
rect 12936 11872 13076 11928
rect 5012 11844 5292 11872
rect 5992 11844 6048 11872
rect 6496 11844 6580 11872
rect 7756 11844 8092 11872
rect 8148 11844 8904 11872
rect 8988 11844 9156 11872
rect 9212 11844 9380 11872
rect 9492 11844 9520 11872
rect 11284 11844 11340 11872
rect 11452 11844 11536 11872
rect 3948 11816 4116 11844
rect 1176 11760 1540 11816
rect 1624 11788 1792 11816
rect 2268 11788 2324 11816
rect 3388 11788 3612 11816
rect 3920 11788 4116 11816
rect 4200 11816 4564 11844
rect 5096 11816 5376 11844
rect 5992 11816 6020 11844
rect 6384 11816 6496 11844
rect 4200 11788 4536 11816
rect 5180 11788 5488 11816
rect 6272 11788 6412 11816
rect 7728 11788 8064 11844
rect 8148 11816 8876 11844
rect 8932 11816 9016 11844
rect 9128 11816 9212 11844
rect 9240 11816 9408 11844
rect 1624 11760 1820 11788
rect 2296 11760 2380 11788
rect 3332 11760 3416 11788
rect 3472 11760 3612 11788
rect 3892 11760 4088 11788
rect 4172 11760 4536 11788
rect 5264 11760 5684 11788
rect 6076 11760 6300 11788
rect 7700 11760 8036 11788
rect 8120 11760 8848 11816
rect 8904 11788 8960 11816
rect 9184 11788 9240 11816
rect 8904 11760 8932 11788
rect 1204 11704 1568 11760
rect 1652 11732 1820 11760
rect 2352 11732 2408 11760
rect 3304 11732 3388 11760
rect 3472 11732 3668 11760
rect 3864 11732 4060 11760
rect 4172 11732 4508 11760
rect 5404 11732 6188 11760
rect 7672 11732 8036 11760
rect 8092 11732 8820 11760
rect 1652 11704 1848 11732
rect 2380 11704 2464 11732
rect 3248 11704 3332 11732
rect 3472 11704 3724 11732
rect 3808 11704 4060 11732
rect 4144 11704 4508 11732
rect 5628 11704 5964 11732
rect 7672 11704 8008 11732
rect 1232 11648 1596 11704
rect 1680 11676 1876 11704
rect 2436 11676 2520 11704
rect 3192 11676 3304 11704
rect 3472 11676 4032 11704
rect 1260 11620 1624 11648
rect 1708 11620 1904 11676
rect 2492 11648 2604 11676
rect 3136 11648 3248 11676
rect 3500 11648 4032 11676
rect 4116 11676 4508 11704
rect 4116 11648 4480 11676
rect 7644 11648 7980 11704
rect 8064 11676 8820 11732
rect 8036 11648 8820 11676
rect 2548 11620 2688 11648
rect 3024 11620 3164 11648
rect 3500 11620 4004 11648
rect 4088 11620 4480 11648
rect 7616 11620 7952 11648
rect 8036 11620 8288 11648
rect 1260 11592 1652 11620
rect 1736 11592 1932 11620
rect 2632 11592 3080 11620
rect 3500 11592 3976 11620
rect 4088 11592 4452 11620
rect 1288 11564 1652 11592
rect 1764 11564 1960 11592
rect 2772 11564 2968 11592
rect 1288 11536 1680 11564
rect 1792 11536 1988 11564
rect 2800 11536 2968 11564
rect 3500 11536 3948 11592
rect 4060 11564 4424 11592
rect 7588 11564 7924 11620
rect 8092 11592 8260 11620
rect 8148 11564 8260 11592
rect 4032 11536 4424 11564
rect 7560 11536 7896 11564
rect 8204 11536 8232 11564
rect 8428 11536 8820 11648
rect 8876 11732 8932 11760
rect 9212 11760 9240 11788
rect 9268 11788 9436 11816
rect 9520 11788 9548 11844
rect 11312 11816 11396 11844
rect 11480 11816 11564 11844
rect 12908 11816 13104 11872
rect 11340 11788 11424 11816
rect 11508 11788 11592 11816
rect 9268 11760 9464 11788
rect 11368 11760 11452 11788
rect 11536 11760 11620 11788
rect 12880 11760 13132 11816
rect 9212 11732 9268 11760
rect 8876 11648 8904 11732
rect 9240 11648 9268 11732
rect 8876 11620 8932 11648
rect 8904 11592 8932 11620
rect 9212 11620 9268 11648
rect 9296 11704 9492 11760
rect 11424 11732 11508 11760
rect 11564 11732 11648 11760
rect 12880 11732 13160 11760
rect 11452 11704 11536 11732
rect 11592 11704 11676 11732
rect 12880 11704 13188 11732
rect 9296 11676 9520 11704
rect 11480 11676 11564 11704
rect 11620 11676 11704 11704
rect 12880 11676 13216 11704
rect 9296 11648 9548 11676
rect 11508 11648 11592 11676
rect 11648 11648 11760 11676
rect 9296 11620 9576 11648
rect 11564 11620 11648 11648
rect 11676 11620 11788 11648
rect 12880 11620 13160 11676
rect 13188 11648 13216 11676
rect 13188 11620 13244 11648
rect 9212 11592 9240 11620
rect 8904 11564 8960 11592
rect 9184 11564 9240 11592
rect 9296 11592 9604 11620
rect 11592 11592 11676 11620
rect 11732 11592 11816 11620
rect 9296 11564 9632 11592
rect 11620 11564 11704 11592
rect 11760 11564 11816 11592
rect 8932 11536 8988 11564
rect 9156 11536 9212 11564
rect 9268 11536 9660 11564
rect 11648 11536 11732 11564
rect 12880 11536 13188 11620
rect 13216 11592 13244 11620
rect 13216 11564 13272 11592
rect 1316 11508 1708 11536
rect 1820 11508 2016 11536
rect 1344 11480 1736 11508
rect 1820 11480 2072 11508
rect 2800 11480 2996 11536
rect 1344 11452 1764 11480
rect 1848 11452 2100 11480
rect 2828 11452 2996 11480
rect 3528 11508 3920 11536
rect 4004 11508 4396 11536
rect 3528 11480 3892 11508
rect 3976 11480 4396 11508
rect 7532 11508 7896 11536
rect 7532 11480 7868 11508
rect 3528 11452 3864 11480
rect 3976 11452 4368 11480
rect 7504 11452 7840 11480
rect 1372 11424 1792 11452
rect 1876 11424 2128 11452
rect 1400 11396 1792 11424
rect 1904 11396 2184 11424
rect 2828 11396 3024 11452
rect 3528 11424 3836 11452
rect 3948 11424 4340 11452
rect 3528 11396 3808 11424
rect 3920 11396 4340 11424
rect 7476 11424 7840 11452
rect 8456 11424 8792 11536
rect 8960 11508 9184 11536
rect 9268 11508 9716 11536
rect 11676 11508 11760 11536
rect 12740 11508 13188 11536
rect 9044 11480 9100 11508
rect 9268 11480 9744 11508
rect 11732 11480 11816 11508
rect 12684 11480 13188 11508
rect 7476 11396 7812 11424
rect 1400 11368 1848 11396
rect 1960 11368 2212 11396
rect 2828 11368 3052 11396
rect 3500 11368 3780 11396
rect 3892 11368 4312 11396
rect 7448 11368 7784 11396
rect 1428 11340 1876 11368
rect 1988 11340 2268 11368
rect 2800 11340 3052 11368
rect 3444 11340 3724 11368
rect 3864 11340 4284 11368
rect 7420 11340 7784 11368
rect 8484 11368 8792 11424
rect 9268 11452 9828 11480
rect 11760 11452 11844 11480
rect 12656 11452 12880 11480
rect 12908 11452 13188 11480
rect 13244 11536 13272 11564
rect 13244 11452 13300 11536
rect 9268 11424 9968 11452
rect 11788 11424 11872 11452
rect 12628 11424 12796 11452
rect 9268 11396 9688 11424
rect 9772 11396 10108 11424
rect 11816 11396 11900 11424
rect 9212 11368 9688 11396
rect 9856 11368 10276 11396
rect 11844 11368 11928 11396
rect 12628 11368 12740 11424
rect 12936 11396 13188 11452
rect 12908 11368 13188 11396
rect 1456 11312 1904 11340
rect 2016 11312 2324 11340
rect 1484 11284 1932 11312
rect 2044 11284 2380 11312
rect 2800 11284 3080 11340
rect 3388 11312 3696 11340
rect 3808 11312 4256 11340
rect 7420 11312 7756 11340
rect 8372 11312 8400 11340
rect 3332 11284 3668 11312
rect 3780 11284 4256 11312
rect 7392 11284 7756 11312
rect 8288 11284 8428 11312
rect 8484 11284 8764 11368
rect 9156 11340 9688 11368
rect 10024 11340 10416 11368
rect 11872 11340 11928 11368
rect 9100 11312 9548 11340
rect 10192 11312 10584 11340
rect 12656 11312 12740 11368
rect 9016 11284 9408 11312
rect 10248 11284 10752 11312
rect 12684 11284 12740 11312
rect 12796 11340 12852 11368
rect 12964 11340 13188 11368
rect 13272 11424 13300 11452
rect 1484 11256 1960 11284
rect 2100 11256 2464 11284
rect 2772 11256 3108 11284
rect 3248 11256 3612 11284
rect 3752 11256 4228 11284
rect 7392 11256 7728 11284
rect 8176 11256 8288 11284
rect 8372 11256 8456 11284
rect 8512 11256 8736 11284
rect 8904 11256 9240 11284
rect 9828 11256 10080 11284
rect 10276 11256 10388 11284
rect 10528 11256 10892 11284
rect 1512 11228 2016 11256
rect 2156 11228 2548 11256
rect 2716 11228 3108 11256
rect 3164 11228 3584 11256
rect 3724 11228 4200 11256
rect 7364 11228 7700 11256
rect 8092 11228 8204 11256
rect 8400 11228 9100 11256
rect 9688 11228 10108 11256
rect 1540 11200 2044 11228
rect 2184 11200 3528 11228
rect 3668 11200 4172 11228
rect 7336 11200 7700 11228
rect 8008 11200 8092 11228
rect 8400 11200 8960 11228
rect 9576 11200 10136 11228
rect 10304 11200 10416 11256
rect 10696 11228 11060 11256
rect 12684 11228 12768 11284
rect 12796 11256 12824 11340
rect 12992 11312 13160 11340
rect 13020 11284 13160 11312
rect 10864 11200 11200 11228
rect 1568 11172 2100 11200
rect 2240 11172 3472 11200
rect 3640 11172 4144 11200
rect 7336 11172 7672 11200
rect 1596 11144 2128 11172
rect 2324 11144 3416 11172
rect 3584 11144 4116 11172
rect 7308 11144 7644 11172
rect 1624 11116 2184 11144
rect 2380 11116 3332 11144
rect 3528 11116 4088 11144
rect 7280 11116 7644 11144
rect 1652 11088 2240 11116
rect 2464 11088 3248 11116
rect 3472 11088 4060 11116
rect 7280 11088 7616 11116
rect 7980 11088 8008 11200
rect 8400 11144 8904 11200
rect 9492 11172 9912 11200
rect 10024 11172 10136 11200
rect 9380 11144 9828 11172
rect 8232 11116 8372 11144
rect 8148 11088 8232 11116
rect 1708 11060 2324 11088
rect 2576 11060 3136 11088
rect 3416 11060 4032 11088
rect 5628 11060 6272 11088
rect 7252 11060 7616 11088
rect 1736 11032 2380 11060
rect 3332 11032 3976 11060
rect 5488 11032 6412 11060
rect 7224 11032 7588 11060
rect 1764 11004 2492 11032
rect 3248 11004 3948 11032
rect 5376 11004 5656 11032
rect 6244 11004 6524 11032
rect 7224 11004 7560 11032
rect 1792 10976 2604 11004
rect 3108 10976 3920 11004
rect 5320 10976 5516 11004
rect 6384 10976 6636 11004
rect 7196 10976 7560 11004
rect 8008 10976 8036 11088
rect 8148 11004 8176 11088
rect 8344 11032 8372 11116
rect 8428 11116 8904 11144
rect 9296 11116 9828 11144
rect 10024 11144 10164 11172
rect 10332 11144 10444 11200
rect 11032 11172 11368 11200
rect 11200 11144 11508 11172
rect 12712 11144 12796 11228
rect 12824 11172 12852 11256
rect 13048 11228 13132 11284
rect 13076 11200 13160 11228
rect 13272 11200 13328 11424
rect 13104 11172 13188 11200
rect 13244 11172 13328 11200
rect 8428 11088 8932 11116
rect 9212 11088 9800 11116
rect 10024 11088 10192 11144
rect 10332 11116 10472 11144
rect 11368 11116 11620 11144
rect 10360 11088 10472 11116
rect 11508 11088 11676 11116
rect 12740 11088 12824 11144
rect 12852 11088 12880 11172
rect 13104 11144 13300 11172
rect 13132 11116 13300 11144
rect 13188 11088 13272 11116
rect 8428 11060 9072 11088
rect 8428 11032 9100 11060
rect 9184 11032 9772 11088
rect 10052 11060 10220 11088
rect 10024 11032 10220 11060
rect 10360 11032 10500 11088
rect 11620 11060 11676 11088
rect 1848 10948 3864 10976
rect 5264 10948 5432 10976
rect 6496 10948 6720 10976
rect 7168 10948 7532 10976
rect 1876 10920 3836 10948
rect 5236 10920 5348 10948
rect 6580 10920 6776 10948
rect 7168 10920 7504 10948
rect 1932 10892 3780 10920
rect 5236 10892 5320 10920
rect 6664 10892 6860 10920
rect 7140 10892 7504 10920
rect 1988 10864 3752 10892
rect 5264 10864 5376 10892
rect 6748 10864 6916 10892
rect 7140 10864 7476 10892
rect 8036 10864 8064 10976
rect 8176 10892 8204 11004
rect 8372 10920 8400 11032
rect 8456 10920 9100 11032
rect 9156 11004 9324 11032
rect 9464 11004 9744 11032
rect 9968 11004 10248 11032
rect 9156 10976 9268 11004
rect 9520 10976 9744 11004
rect 9856 10976 10248 11004
rect 9156 10948 9240 10976
rect 2016 10836 3696 10864
rect 5292 10836 5488 10864
rect 6832 10836 6972 10864
rect 7112 10836 7476 10864
rect 2072 10808 3640 10836
rect 5320 10808 5656 10836
rect 6888 10808 7028 10836
rect 7084 10808 7448 10836
rect 2156 10780 3584 10808
rect 5236 10780 5880 10808
rect 6944 10780 7420 10808
rect 2212 10752 3500 10780
rect 5152 10752 6076 10780
rect 7000 10752 7420 10780
rect 8064 10752 8092 10864
rect 8204 10780 8232 10892
rect 8400 10808 8428 10920
rect 8484 10836 9128 10920
rect 9156 10892 9268 10948
rect 9576 10920 10276 10976
rect 10388 10920 10528 11032
rect 12768 11004 12852 11088
rect 12880 11004 12908 11088
rect 12796 10948 12880 11004
rect 12824 10920 12880 10948
rect 12908 10920 12936 11004
rect 9548 10892 10304 10920
rect 9156 10864 9296 10892
rect 9464 10864 9744 10892
rect 2296 10724 3416 10752
rect 5096 10724 6216 10752
rect 7028 10724 7392 10752
rect 2380 10696 3332 10724
rect 5040 10696 6328 10724
rect 7028 10696 7364 10724
rect 2520 10668 3220 10696
rect 4984 10668 6412 10696
rect 7000 10668 7364 10696
rect 8092 10668 8120 10752
rect 8232 10668 8260 10780
rect 8428 10696 8456 10808
rect 8512 10780 9128 10836
rect 9184 10836 9296 10864
rect 9380 10836 9604 10864
rect 8512 10724 9156 10780
rect 9184 10724 9632 10836
rect 9688 10780 9744 10864
rect 9800 10864 10304 10892
rect 9800 10836 10192 10864
rect 10248 10836 10304 10864
rect 10388 10836 10556 10920
rect 10752 10836 11228 10864
rect 12404 10836 12768 10920
rect 12824 10864 12908 10920
rect 12936 10864 12964 10920
rect 12852 10836 12964 10864
rect 15008 10836 15092 11088
rect 15288 11004 15372 11088
rect 15260 10920 15344 11004
rect 15484 10976 15568 11088
rect 15680 10976 15820 11088
rect 15988 11004 16072 11088
rect 16296 11060 16492 11088
rect 16660 11060 16940 11088
rect 16268 11032 16520 11060
rect 15456 10948 15568 10976
rect 15232 10836 15316 10920
rect 15456 10836 15540 10948
rect 15652 10920 15820 10976
rect 15652 10836 15736 10920
rect 9800 10808 10080 10836
rect 10192 10808 10332 10836
rect 10388 10808 11396 10836
rect 9828 10780 9968 10808
rect 10080 10780 10248 10808
rect 10388 10780 10808 10808
rect 11200 10780 11480 10808
rect 9688 10752 9772 10780
rect 9828 10752 9856 10780
rect 9968 10752 10108 10780
rect 10332 10752 10612 10780
rect 11368 10752 11452 10780
rect 9716 10724 9744 10752
rect 9856 10724 9996 10752
rect 10360 10724 10472 10752
rect 2716 10640 2996 10668
rect 4928 10640 6524 10668
rect 4872 10612 6580 10640
rect 6972 10612 7336 10668
rect 8092 10640 8148 10668
rect 4816 10584 6664 10612
rect 6944 10584 7364 10612
rect 4788 10556 6720 10584
rect 6916 10556 7392 10584
rect 8120 10556 8148 10640
rect 8260 10556 8288 10668
rect 8456 10584 8484 10696
rect 8540 10612 9156 10724
rect 9212 10696 9632 10724
rect 9744 10696 9884 10724
rect 10192 10696 10332 10724
rect 9212 10668 9520 10696
rect 9632 10668 9772 10696
rect 10080 10668 10332 10696
rect 10360 10696 10416 10724
rect 9212 10640 9408 10668
rect 9520 10640 9660 10668
rect 9968 10640 10220 10668
rect 10360 10640 10444 10696
rect 9212 10612 9296 10640
rect 9408 10612 9548 10640
rect 9856 10612 10108 10640
rect 10248 10612 10360 10640
rect 4732 10528 6776 10556
rect 6916 10528 7280 10556
rect 7336 10528 7420 10556
rect 4704 10500 5628 10528
rect 6188 10500 6832 10528
rect 6888 10500 7252 10528
rect 7364 10500 7448 10528
rect 4676 10472 5488 10500
rect 6328 10472 7224 10500
rect 7392 10472 7476 10500
rect 4620 10444 5404 10472
rect 6412 10444 7224 10472
rect 7420 10444 7504 10472
rect 8148 10444 8176 10556
rect 8288 10444 8316 10556
rect 8484 10472 8512 10584
rect 8568 10500 9184 10612
rect 9240 10584 9436 10612
rect 9744 10584 9996 10612
rect 10136 10584 10360 10612
rect 10388 10584 10444 10640
rect 12404 10612 12432 10836
rect 12600 10780 12656 10808
rect 12572 10752 12684 10780
rect 12712 10752 12740 10836
rect 12852 10808 12936 10836
rect 12964 10808 12992 10836
rect 12572 10724 12600 10752
rect 12684 10724 12740 10752
rect 12880 10752 12992 10808
rect 12880 10724 13020 10752
rect 12544 10696 12572 10724
rect 12712 10696 12768 10724
rect 12516 10668 12572 10696
rect 12740 10668 12824 10696
rect 12908 10668 13020 10724
rect 13188 10696 13384 10724
rect 13132 10668 13440 10696
rect 13496 10668 13636 10696
rect 12488 10640 12544 10668
rect 12684 10640 12740 10668
rect 12796 10640 12852 10668
rect 12936 10640 13048 10668
rect 13104 10640 13692 10668
rect 12488 10612 12516 10640
rect 12656 10612 12712 10640
rect 12852 10612 12908 10640
rect 12936 10612 13524 10640
rect 13636 10612 13720 10640
rect 12432 10584 12488 10612
rect 12656 10584 12684 10612
rect 12880 10584 13468 10612
rect 9240 10556 9324 10584
rect 9632 10556 9912 10584
rect 10024 10556 10304 10584
rect 9520 10528 9800 10556
rect 9940 10528 10192 10556
rect 10332 10528 10360 10556
rect 10388 10528 10472 10584
rect 12432 10556 12460 10584
rect 12628 10556 12656 10584
rect 12936 10556 13412 10584
rect 11480 10528 11592 10556
rect 12404 10528 12460 10556
rect 12600 10528 12628 10556
rect 12964 10528 13356 10556
rect 9408 10500 9688 10528
rect 9828 10500 10080 10528
rect 10220 10500 10388 10528
rect 8596 10472 9100 10500
rect 9324 10472 9576 10500
rect 9716 10472 9968 10500
rect 10108 10472 10360 10500
rect 10416 10472 10472 10528
rect 11452 10500 11620 10528
rect 12404 10500 12432 10528
rect 12572 10500 12628 10528
rect 12992 10500 13300 10528
rect 13664 10500 13720 10612
rect 14980 10528 15064 10836
rect 15204 10752 15288 10836
rect 15176 10696 15260 10752
rect 15428 10696 15512 10836
rect 15624 10696 15708 10836
rect 15176 10668 15232 10696
rect 15148 10612 15232 10668
rect 15120 10528 15204 10612
rect 15400 10584 15484 10696
rect 15596 10584 15680 10696
rect 15372 10556 15484 10584
rect 15568 10556 15680 10584
rect 10612 10472 11060 10500
rect 11424 10472 11508 10500
rect 11564 10472 11648 10500
rect 12376 10472 12404 10500
rect 12572 10472 12600 10500
rect 12768 10472 13160 10500
rect 13636 10472 13692 10500
rect 14980 10472 15036 10528
rect 4592 10416 5320 10444
rect 5684 10416 6132 10444
rect 6496 10416 7196 10444
rect 7448 10416 7532 10444
rect 4564 10388 5236 10416
rect 5516 10388 6300 10416
rect 6580 10388 7168 10416
rect 7476 10388 7560 10416
rect 4536 10360 5180 10388
rect 5432 10360 6384 10388
rect 6636 10360 7168 10388
rect 7504 10360 7588 10388
rect 4508 10332 5124 10360
rect 5348 10332 6468 10360
rect 6692 10332 7140 10360
rect 7532 10332 7616 10360
rect 8176 10332 8204 10444
rect 8316 10332 8344 10444
rect 8512 10360 8540 10472
rect 8596 10388 8988 10472
rect 4480 10304 5068 10332
rect 5264 10304 6552 10332
rect 6748 10304 7168 10332
rect 7560 10304 7616 10332
rect 4452 10276 5040 10304
rect 5208 10276 6608 10304
rect 6748 10276 7196 10304
rect 7560 10276 7644 10304
rect 4424 10248 4984 10276
rect 5152 10248 6664 10276
rect 6720 10248 7224 10276
rect 7588 10248 7672 10276
rect 4396 10220 4956 10248
rect 5096 10220 5572 10248
rect 5684 10220 6104 10248
rect 6244 10220 7252 10248
rect 4368 10192 4900 10220
rect 5068 10192 5488 10220
rect 4340 10164 4872 10192
rect 5012 10164 5404 10192
rect 5712 10164 5880 10220
rect 4312 10136 4844 10164
rect 4984 10136 5348 10164
rect 5740 10136 5880 10164
rect 4284 10108 4788 10136
rect 4928 10108 5264 10136
rect 4284 10080 4760 10108
rect 4900 10080 5236 10108
rect 5768 10080 5880 10136
rect 4256 10052 4732 10080
rect 4872 10052 5180 10080
rect 4228 10024 4704 10052
rect 4844 10024 5124 10052
rect 4200 9996 4676 10024
rect 4816 9996 5096 10024
rect 4200 9968 4648 9996
rect 4788 9968 5040 9996
rect 4172 9940 4620 9968
rect 4760 9940 5012 9968
rect 4144 9912 4620 9940
rect 4732 9912 4984 9940
rect 4144 9884 4592 9912
rect 4704 9884 4956 9912
rect 5796 9884 5880 10080
rect 4116 9856 4564 9884
rect 4676 9856 4928 9884
rect 4116 9828 4536 9856
rect 4648 9828 4900 9856
rect 4088 9800 4536 9828
rect 4620 9800 4872 9828
rect 4088 9772 4508 9800
rect 4620 9772 4844 9800
rect 5824 9772 5880 9884
rect 5908 10192 6076 10220
rect 6328 10192 7280 10220
rect 7616 10192 7700 10248
rect 8204 10220 8232 10332
rect 8344 10248 8372 10332
rect 8540 10248 8568 10360
rect 8624 10304 8988 10388
rect 9072 10444 9100 10472
rect 9212 10444 9464 10472
rect 9604 10444 9856 10472
rect 9996 10444 10248 10472
rect 10416 10444 11060 10472
rect 11396 10444 11480 10472
rect 11592 10444 11676 10472
rect 12348 10444 12376 10472
rect 12488 10444 12964 10472
rect 13608 10444 13692 10472
rect 9072 10416 9352 10444
rect 9492 10416 9744 10444
rect 9884 10416 10136 10444
rect 10276 10416 10388 10444
rect 10416 10416 10668 10444
rect 11004 10416 11032 10444
rect 9072 10388 9240 10416
rect 9380 10388 9632 10416
rect 9772 10388 10024 10416
rect 10164 10388 10388 10416
rect 10444 10388 10500 10416
rect 11396 10388 11452 10444
rect 11620 10416 11704 10444
rect 12320 10416 12740 10444
rect 13552 10416 13664 10444
rect 11648 10388 11732 10416
rect 12292 10388 12460 10416
rect 13496 10388 13636 10416
rect 9072 10360 9128 10388
rect 9268 10360 9520 10388
rect 9660 10360 9912 10388
rect 10052 10360 10304 10388
rect 10556 10360 10612 10388
rect 11396 10360 11480 10388
rect 11676 10360 11760 10388
rect 12236 10360 12376 10388
rect 13412 10360 13580 10388
rect 9100 10332 9128 10360
rect 9156 10332 9408 10360
rect 9548 10332 9800 10360
rect 9940 10332 10192 10360
rect 10444 10332 10724 10360
rect 11424 10332 11480 10360
rect 11704 10332 11788 10360
rect 12236 10332 12320 10360
rect 13300 10332 13524 10360
rect 9100 10304 9296 10332
rect 9436 10304 9688 10332
rect 9828 10304 10080 10332
rect 10388 10304 10472 10332
rect 10696 10304 10752 10332
rect 11424 10304 11508 10332
rect 11732 10304 11816 10332
rect 8652 10276 8960 10304
rect 9100 10276 9184 10304
rect 9324 10276 9576 10304
rect 9716 10276 9968 10304
rect 10360 10276 10416 10304
rect 10724 10276 10780 10304
rect 11396 10276 11536 10304
rect 11760 10276 11816 10304
rect 8652 10248 8932 10276
rect 9044 10248 9128 10276
rect 9212 10248 9464 10276
rect 9604 10248 9884 10276
rect 10332 10248 10388 10276
rect 10780 10248 10808 10276
rect 8344 10220 8400 10248
rect 5908 10164 6048 10192
rect 6412 10164 7308 10192
rect 7644 10164 7728 10192
rect 5908 10108 6020 10164
rect 6468 10136 7336 10164
rect 7672 10136 7728 10164
rect 6552 10108 7364 10136
rect 7672 10108 7756 10136
rect 8232 10108 8260 10220
rect 8372 10136 8400 10220
rect 8568 10164 8596 10248
rect 8652 10220 8904 10248
rect 8988 10220 9100 10248
rect 8652 10192 8848 10220
rect 8960 10192 9100 10220
rect 8484 10136 8596 10164
rect 8680 10164 8820 10192
rect 8904 10164 8988 10192
rect 9044 10164 9100 10192
rect 8680 10136 8792 10164
rect 8876 10136 8960 10164
rect 9072 10136 9100 10164
rect 9128 10220 9380 10248
rect 9492 10220 9772 10248
rect 10304 10220 10360 10248
rect 10780 10220 10836 10248
rect 11396 10220 11452 10276
rect 11480 10248 11564 10276
rect 11788 10248 11844 10276
rect 12236 10248 12292 10332
rect 13132 10304 13524 10332
rect 12824 10276 13524 10304
rect 12516 10248 13524 10276
rect 14952 10332 15036 10472
rect 15092 10444 15176 10528
rect 15372 10444 15456 10556
rect 15568 10444 15652 10556
rect 15064 10360 15148 10444
rect 15064 10332 15120 10360
rect 14952 10276 15120 10332
rect 15344 10304 15428 10444
rect 15540 10304 15624 10444
rect 15764 10416 15820 10920
rect 15960 10976 16072 11004
rect 16212 11004 16520 11032
rect 16660 11004 16912 11060
rect 16212 10976 16324 11004
rect 15960 10864 16044 10976
rect 16184 10948 16296 10976
rect 16184 10864 16268 10948
rect 15932 10836 16044 10864
rect 16156 10836 16268 10864
rect 16436 10920 16548 11004
rect 16660 10976 16744 11004
rect 17052 10976 17192 11088
rect 17360 11004 17444 11088
rect 17528 11060 17836 11088
rect 18088 11060 18368 11088
rect 17500 11004 17808 11060
rect 18088 11004 18340 11060
rect 16632 10948 16744 10976
rect 15932 10724 16016 10836
rect 16156 10724 16240 10836
rect 16436 10808 16520 10920
rect 16632 10836 16716 10948
rect 17024 10920 17192 10976
rect 17024 10836 17108 10920
rect 16408 10780 16492 10808
rect 16604 10724 16688 10836
rect 15904 10612 15988 10724
rect 15876 10584 15988 10612
rect 16128 10584 16212 10724
rect 16604 10696 16828 10724
rect 16996 10696 17080 10836
rect 16576 10640 16828 10696
rect 16576 10584 16660 10640
rect 16968 10584 17052 10696
rect 15876 10444 15960 10584
rect 16100 10472 16184 10584
rect 16548 10556 16660 10584
rect 16940 10556 17052 10584
rect 16072 10444 16184 10472
rect 16352 10528 16464 10556
rect 15848 10416 15932 10444
rect 15764 10332 15932 10416
rect 16072 10360 16156 10444
rect 16352 10416 16436 10528
rect 16548 10444 16632 10556
rect 16940 10444 17024 10556
rect 16324 10388 16436 10416
rect 16324 10360 16408 10388
rect 16072 10332 16184 10360
rect 16296 10332 16408 10360
rect 16520 10332 16604 10444
rect 14952 10248 15092 10276
rect 15316 10248 15400 10304
rect 15512 10248 15596 10304
rect 15764 10248 15904 10332
rect 16072 10304 16380 10332
rect 16520 10304 16772 10332
rect 16912 10304 16996 10444
rect 17136 10416 17192 10920
rect 17332 10976 17444 11004
rect 17332 10864 17416 10976
rect 17612 10920 17696 11004
rect 18088 10976 18172 11004
rect 18452 10976 18536 11088
rect 18732 11060 18816 11088
rect 18984 11060 19180 11088
rect 19460 11060 19656 11088
rect 19908 11060 20104 11088
rect 18060 10948 18172 10976
rect 17304 10836 17416 10864
rect 17304 10724 17388 10836
rect 17584 10808 17668 10920
rect 18060 10836 18144 10948
rect 18424 10836 18508 10976
rect 18704 10920 18788 11060
rect 18956 11032 19208 11060
rect 19432 11032 19684 11060
rect 19880 11032 20132 11060
rect 18928 11004 19236 11032
rect 18900 10976 19012 11004
rect 19124 10976 19236 11004
rect 19376 11004 19684 11032
rect 19824 11004 20132 11032
rect 19376 10976 19488 11004
rect 18900 10920 18984 10976
rect 17556 10780 17668 10808
rect 17276 10612 17360 10724
rect 17556 10668 17640 10780
rect 18032 10724 18116 10836
rect 18396 10724 18480 10836
rect 18676 10808 18760 10920
rect 18872 10808 18956 10920
rect 19152 10892 19236 10976
rect 19348 10948 19460 10976
rect 19124 10836 19208 10892
rect 19348 10864 19432 10948
rect 19320 10836 19432 10864
rect 19600 10920 19712 11004
rect 19824 10976 19936 11004
rect 19796 10948 19908 10976
rect 18032 10696 18256 10724
rect 17248 10584 17360 10612
rect 17528 10640 17640 10668
rect 18004 10640 18256 10696
rect 18368 10696 18480 10724
rect 18648 10780 18760 10808
rect 18844 10780 18956 10808
rect 17248 10444 17332 10584
rect 17528 10528 17612 10640
rect 18004 10584 18088 10640
rect 18368 10584 18452 10696
rect 18648 10668 18732 10780
rect 18844 10752 18984 10780
rect 18872 10724 19012 10752
rect 19320 10724 19404 10836
rect 19600 10808 19684 10920
rect 19796 10864 19880 10948
rect 19768 10836 19880 10864
rect 20048 10920 20160 11004
rect 19572 10780 19656 10808
rect 19768 10724 19852 10836
rect 20048 10808 20132 10920
rect 18900 10696 19040 10724
rect 18928 10668 19068 10696
rect 17976 10556 18088 10584
rect 17220 10416 17304 10444
rect 17136 10332 17304 10416
rect 17500 10388 17584 10528
rect 17976 10444 18060 10556
rect 18340 10444 18424 10584
rect 18620 10528 18704 10668
rect 18956 10640 19096 10668
rect 18984 10612 19124 10640
rect 19012 10584 19152 10612
rect 19292 10584 19376 10724
rect 19740 10584 19824 10724
rect 20020 10668 20104 10808
rect 19040 10556 19152 10584
rect 16100 10276 16352 10304
rect 16128 10248 16324 10276
rect 16492 10248 16772 10304
rect 16884 10248 16968 10304
rect 17136 10248 17276 10332
rect 17472 10276 17556 10388
rect 17948 10304 18032 10444
rect 18312 10360 18396 10444
rect 18592 10416 18676 10528
rect 18788 10416 18872 10528
rect 19068 10500 19152 10556
rect 18564 10388 18676 10416
rect 18564 10360 18648 10388
rect 18312 10332 18424 10360
rect 18536 10332 18648 10360
rect 18760 10332 18872 10416
rect 19040 10472 19152 10500
rect 19264 10472 19348 10584
rect 19040 10388 19124 10472
rect 19012 10360 19124 10388
rect 19236 10444 19348 10472
rect 19516 10528 19628 10556
rect 19236 10360 19320 10444
rect 19516 10416 19600 10528
rect 19712 10472 19796 10584
rect 19992 10556 20076 10668
rect 19488 10388 19600 10416
rect 19684 10444 19796 10472
rect 19964 10528 20076 10556
rect 19488 10360 19572 10388
rect 18984 10332 19096 10360
rect 18312 10304 18620 10332
rect 18788 10304 19096 10332
rect 19236 10332 19348 10360
rect 19460 10332 19572 10360
rect 19684 10360 19768 10444
rect 19964 10416 20048 10528
rect 19936 10388 20048 10416
rect 19936 10360 20020 10388
rect 19684 10332 19796 10360
rect 19908 10332 20020 10360
rect 19236 10304 19544 10332
rect 19684 10304 19992 10332
rect 17444 10248 17556 10276
rect 17920 10248 18004 10304
rect 18340 10276 18592 10304
rect 18788 10276 19040 10304
rect 19264 10276 19516 10304
rect 19712 10276 19964 10304
rect 18368 10248 18564 10276
rect 18816 10248 19012 10276
rect 19292 10248 19488 10276
rect 19740 10248 19936 10276
rect 11508 10220 11592 10248
rect 11788 10220 11872 10248
rect 9128 10192 9268 10220
rect 9380 10192 9660 10220
rect 9828 10192 9912 10220
rect 9996 10192 10052 10220
rect 10304 10192 10332 10220
rect 10808 10192 10864 10220
rect 11396 10192 11480 10220
rect 11508 10192 11620 10220
rect 11816 10192 11900 10220
rect 12264 10192 12320 10248
rect 12488 10220 12740 10248
rect 13076 10220 13524 10248
rect 12460 10192 12544 10220
rect 13048 10192 13524 10220
rect 9128 10164 9156 10192
rect 9296 10164 9548 10192
rect 9716 10164 9800 10192
rect 10052 10164 10136 10192
rect 9128 10136 9436 10164
rect 9632 10136 9688 10164
rect 9968 10136 10136 10164
rect 10276 10164 10332 10192
rect 8400 10108 8484 10136
rect 8680 10108 8764 10136
rect 8848 10108 8932 10136
rect 5908 10052 5992 10108
rect 6580 10080 7000 10108
rect 7056 10080 7392 10108
rect 7700 10080 7756 10108
rect 6608 10052 6972 10080
rect 7084 10052 7420 10080
rect 7700 10052 7784 10080
rect 5908 9772 5964 10052
rect 6580 10024 6972 10052
rect 7112 10024 7448 10052
rect 7728 10024 7784 10052
rect 8260 10024 8288 10108
rect 8680 10052 8736 10108
rect 8820 10080 8904 10108
rect 8792 10052 8876 10080
rect 9072 10052 9128 10136
rect 8652 10024 8680 10052
rect 8764 10024 8848 10052
rect 9100 10024 9128 10052
rect 9156 10108 9324 10136
rect 9576 10108 9632 10136
rect 9856 10108 9968 10136
rect 10108 10108 10164 10136
rect 9156 10080 9212 10108
rect 9576 10080 9604 10108
rect 9716 10080 9856 10108
rect 10052 10080 10164 10108
rect 9156 10024 9184 10080
rect 9548 10052 9576 10080
rect 9604 10052 9716 10080
rect 9940 10052 10052 10080
rect 10136 10052 10164 10080
rect 9492 10024 9604 10052
rect 9800 10024 9940 10052
rect 6580 9996 7000 10024
rect 7140 9996 7476 10024
rect 7728 9996 7812 10024
rect 6552 9968 7028 9996
rect 7168 9968 7504 9996
rect 7756 9968 7812 9996
rect 6524 9940 7056 9968
rect 6524 9912 7084 9940
rect 7196 9912 7532 9968
rect 7756 9940 7840 9968
rect 7784 9912 7840 9940
rect 8288 9940 8316 10024
rect 8624 9996 8652 10024
rect 8736 9996 8820 10024
rect 9072 9996 9212 10024
rect 8568 9968 8624 9996
rect 8708 9968 8792 9996
rect 9044 9968 9128 9996
rect 9184 9968 9212 9996
rect 9520 9968 9548 10024
rect 9688 9996 9800 10024
rect 9576 9968 9688 9996
rect 10164 9968 10192 10052
rect 10276 9968 10304 10164
rect 10836 10136 10864 10192
rect 11424 10164 11508 10192
rect 11536 10164 11620 10192
rect 11844 10164 11928 10192
rect 12264 10164 12348 10192
rect 12432 10164 12516 10192
rect 12992 10164 13496 10192
rect 11452 10136 11648 10164
rect 11872 10136 11956 10164
rect 12292 10136 12488 10164
rect 12908 10136 13216 10164
rect 13272 10136 13412 10164
rect 10836 10108 10892 10136
rect 11508 10108 11564 10136
rect 11592 10108 11676 10136
rect 11900 10108 11984 10136
rect 12320 10108 12432 10136
rect 12656 10108 13188 10136
rect 13300 10108 13328 10136
rect 10864 10052 10892 10108
rect 11592 10080 11704 10108
rect 11928 10080 11984 10108
rect 12348 10080 12432 10108
rect 12628 10080 13160 10108
rect 11536 10052 11732 10080
rect 11956 10052 12012 10080
rect 12292 10052 12376 10080
rect 12432 10052 12460 10080
rect 12600 10052 13160 10080
rect 14784 10052 20076 10108
rect 10836 9996 10892 10052
rect 11508 10024 11760 10052
rect 11956 10024 12040 10052
rect 12236 10024 12348 10052
rect 12432 10024 12516 10052
rect 12572 10024 13104 10052
rect 14756 10024 20076 10052
rect 8540 9940 8596 9968
rect 8680 9940 8764 9968
rect 9016 9940 9100 9968
rect 9184 9940 9240 9968
rect 9492 9940 9576 9968
rect 10276 9940 10332 9968
rect 10836 9940 10864 9996
rect 11508 9968 11788 10024
rect 11116 9940 11172 9968
rect 11480 9940 11816 9968
rect 8288 9912 8344 9940
rect 8512 9912 8568 9940
rect 8652 9912 8736 9940
rect 8988 9912 9072 9940
rect 6496 9884 7112 9912
rect 7224 9884 7560 9912
rect 7784 9884 7868 9912
rect 6468 9856 6860 9884
rect 6888 9856 7140 9884
rect 7252 9856 7588 9884
rect 6468 9828 6832 9856
rect 6916 9828 7168 9856
rect 7280 9828 7588 9856
rect 7812 9828 7868 9884
rect 8624 9884 8708 9912
rect 8960 9884 9072 9912
rect 9184 9912 9296 9940
rect 9184 9884 9324 9912
rect 8624 9856 8680 9884
rect 8932 9856 9100 9884
rect 9184 9856 9352 9884
rect 8596 9828 8680 9856
rect 8904 9828 8988 9856
rect 9016 9828 9100 9856
rect 6440 9800 6804 9828
rect 6944 9800 7196 9828
rect 7280 9800 7616 9828
rect 7812 9800 7896 9828
rect 8596 9800 8652 9828
rect 8904 9800 8960 9828
rect 4060 9716 4480 9772
rect 4592 9744 4816 9772
rect 5796 9744 5964 9772
rect 6412 9772 6804 9800
rect 6972 9772 7196 9800
rect 7308 9772 7644 9800
rect 6412 9744 6776 9772
rect 7000 9744 7224 9772
rect 7336 9744 7644 9772
rect 7840 9772 7896 9800
rect 8568 9772 8624 9800
rect 8876 9772 8960 9800
rect 9044 9772 9100 9828
rect 9212 9828 9380 9856
rect 9520 9828 9548 9912
rect 10192 9828 10220 9940
rect 10304 9912 10332 9940
rect 10808 9912 10836 9940
rect 11060 9912 11144 9940
rect 11452 9912 11844 9940
rect 11984 9912 12040 10024
rect 12180 9996 12292 10024
rect 12404 9996 13020 10024
rect 14756 9996 20048 10024
rect 12152 9968 12264 9996
rect 12348 9968 12908 9996
rect 14728 9968 20048 9996
rect 12096 9940 12236 9968
rect 12292 9940 12460 9968
rect 12544 9940 12880 9968
rect 14728 9940 20020 9968
rect 12068 9912 12432 9940
rect 12516 9912 12824 9940
rect 14728 9912 19992 9940
rect 10332 9884 10360 9912
rect 10780 9884 10836 9912
rect 11004 9884 11088 9912
rect 11452 9884 11900 9912
rect 11928 9884 12376 9912
rect 12516 9884 12796 9912
rect 14700 9884 19992 9912
rect 10332 9856 10388 9884
rect 10752 9856 10808 9884
rect 10920 9856 11004 9884
rect 11452 9856 12348 9884
rect 12516 9856 12740 9884
rect 10360 9828 10416 9856
rect 10724 9828 10780 9856
rect 10836 9828 10948 9856
rect 11508 9828 11788 9856
rect 11872 9828 11956 9856
rect 11984 9828 12292 9856
rect 9212 9800 9436 9828
rect 10388 9800 10472 9828
rect 10668 9800 10864 9828
rect 11564 9800 11788 9828
rect 11956 9800 12320 9828
rect 12488 9800 12712 9856
rect 9212 9772 9464 9800
rect 4564 9716 4788 9744
rect 5712 9716 6104 9744
rect 4032 9688 4452 9716
rect 4564 9688 4760 9716
rect 5600 9688 6216 9716
rect 6384 9688 6748 9744
rect 7028 9716 7252 9744
rect 7336 9716 7672 9744
rect 7840 9716 7924 9772
rect 7056 9688 7252 9716
rect 7364 9688 7672 9716
rect 4032 9660 4424 9688
rect 4536 9660 4760 9688
rect 5544 9660 5740 9688
rect 6076 9660 6272 9688
rect 6356 9660 6720 9688
rect 7056 9660 7280 9688
rect 4004 9632 4424 9660
rect 4508 9632 4732 9660
rect 5488 9632 5656 9660
rect 6160 9632 6720 9660
rect 7084 9632 7308 9660
rect 7392 9632 7700 9688
rect 7868 9660 7924 9716
rect 8540 9744 8624 9772
rect 8848 9744 8932 9772
rect 8540 9688 8596 9744
rect 8848 9716 8960 9744
rect 9044 9716 9128 9772
rect 9212 9744 9240 9772
rect 9296 9744 9492 9772
rect 8512 9660 8596 9688
rect 8820 9688 8960 9716
rect 7868 9632 7952 9660
rect 4004 9576 4396 9632
rect 4508 9604 4704 9632
rect 5432 9604 5572 9632
rect 6244 9604 6692 9632
rect 7112 9604 7308 9632
rect 4480 9576 4704 9604
rect 5376 9576 5516 9604
rect 6300 9576 6664 9604
rect 3976 9520 4368 9576
rect 4480 9548 4676 9576
rect 5348 9548 5460 9576
rect 6272 9548 6664 9576
rect 7112 9548 7336 9604
rect 7420 9576 7728 9632
rect 4452 9520 4676 9548
rect 5320 9520 5432 9548
rect 6272 9520 6636 9548
rect 7112 9520 7364 9548
rect 7448 9520 7756 9576
rect 7896 9548 7952 9632
rect 8512 9604 8568 9660
rect 8820 9632 8876 9688
rect 8904 9632 8960 9688
rect 9072 9660 9128 9716
rect 9240 9660 9268 9744
rect 9352 9716 9520 9744
rect 9380 9688 9520 9716
rect 9548 9688 9576 9800
rect 10192 9716 10220 9800
rect 10444 9772 10780 9800
rect 11592 9772 11788 9800
rect 11928 9772 12376 9800
rect 12460 9772 12684 9800
rect 13468 9772 13888 9800
rect 10528 9744 10696 9772
rect 11172 9744 11284 9772
rect 11648 9744 11844 9772
rect 11928 9744 12152 9772
rect 12180 9744 12656 9772
rect 13384 9744 13468 9772
rect 10444 9716 10612 9744
rect 11144 9716 11284 9744
rect 11676 9716 12124 9744
rect 10164 9688 10192 9716
rect 10360 9688 10528 9716
rect 8484 9576 8568 9604
rect 7896 9520 7980 9548
rect 3948 9436 4340 9520
rect 4452 9492 4648 9520
rect 5292 9492 5376 9520
rect 6244 9492 6608 9520
rect 4424 9436 4676 9492
rect 5264 9464 5348 9492
rect 6216 9464 6608 9492
rect 7084 9492 7364 9520
rect 7084 9464 7392 9492
rect 5236 9436 5320 9464
rect 6216 9436 6636 9464
rect 7056 9436 7392 9464
rect 7476 9464 7784 9520
rect 7476 9436 7812 9464
rect 3948 9408 4312 9436
rect 4424 9408 4704 9436
rect 5208 9408 5292 9436
rect 5768 9408 6048 9436
rect 6188 9408 6692 9436
rect 7028 9408 7392 9436
rect 3920 9352 4312 9408
rect 4396 9380 4704 9408
rect 5180 9380 5264 9408
rect 5684 9380 5936 9408
rect 5964 9380 6132 9408
rect 6160 9380 6804 9408
rect 7000 9380 7420 9408
rect 4396 9352 4732 9380
rect 3920 9296 4284 9352
rect 4396 9324 4760 9352
rect 5152 9324 5236 9380
rect 5628 9352 5740 9380
rect 5572 9324 5656 9352
rect 3892 9268 4284 9296
rect 4368 9296 4788 9324
rect 5124 9296 5208 9324
rect 5544 9296 5656 9324
rect 4368 9268 4816 9296
rect 5124 9268 5180 9296
rect 5516 9268 5656 9296
rect 5796 9296 5908 9380
rect 6076 9324 6524 9380
rect 6552 9352 6804 9380
rect 6972 9352 7140 9380
rect 7196 9352 7420 9380
rect 7504 9380 7812 9436
rect 7924 9380 7980 9520
rect 8484 9380 8540 9576
rect 8792 9520 8848 9632
rect 8904 9576 8988 9632
rect 9072 9604 9156 9660
rect 9240 9632 9296 9660
rect 8932 9520 8988 9576
rect 9100 9576 9156 9604
rect 9268 9576 9296 9632
rect 9408 9576 9520 9688
rect 9576 9632 9604 9688
rect 10136 9660 10164 9688
rect 10248 9660 10416 9688
rect 10108 9632 10332 9660
rect 9604 9604 9632 9632
rect 9996 9604 10220 9632
rect 9632 9576 9688 9604
rect 9856 9576 10108 9604
rect 9100 9520 9184 9576
rect 9268 9548 9380 9576
rect 9408 9548 9548 9576
rect 9604 9548 9968 9576
rect 9268 9520 9856 9548
rect 9912 9520 10192 9548
rect 8764 9436 8820 9520
rect 8932 9492 9016 9520
rect 8960 9436 9016 9492
rect 9128 9464 9184 9520
rect 9296 9492 9604 9520
rect 9828 9492 10248 9520
rect 9296 9464 9324 9492
rect 9772 9464 10304 9492
rect 7504 9352 7840 9380
rect 6580 9324 6804 9352
rect 6916 9324 7084 9352
rect 7140 9324 7420 9352
rect 7532 9324 7840 9352
rect 7924 9324 8008 9380
rect 8484 9352 8568 9380
rect 6048 9296 6496 9324
rect 6608 9296 6832 9324
rect 6860 9296 7028 9324
rect 7084 9296 7448 9324
rect 3892 9156 4256 9268
rect 4368 9240 4620 9268
rect 4676 9240 4900 9268
rect 5096 9240 5180 9268
rect 5488 9240 5684 9268
rect 5796 9240 5936 9296
rect 6048 9268 6468 9296
rect 6580 9268 6972 9296
rect 7028 9268 7448 9296
rect 7532 9296 7868 9324
rect 7532 9268 7896 9296
rect 6020 9240 6468 9268
rect 6552 9240 6916 9268
rect 6972 9240 7448 9268
rect 4368 9212 4704 9240
rect 4760 9212 4984 9240
rect 5096 9212 5152 9240
rect 5460 9212 5516 9240
rect 5544 9212 5712 9240
rect 5796 9212 6440 9240
rect 3864 9128 4256 9156
rect 4340 9184 4788 9212
rect 4844 9184 5152 9212
rect 5432 9184 5488 9212
rect 5572 9184 5796 9212
rect 6020 9184 6440 9212
rect 6524 9212 6860 9240
rect 6916 9212 7084 9240
rect 7196 9212 7448 9240
rect 7560 9240 7924 9268
rect 7952 9240 8008 9324
rect 8512 9296 8568 9352
rect 8792 9324 8848 9436
rect 8960 9380 9044 9436
rect 9128 9408 9212 9464
rect 9296 9436 9352 9464
rect 9744 9436 10360 9464
rect 8988 9352 9044 9380
rect 9156 9380 9212 9408
rect 9324 9380 9352 9436
rect 9716 9408 10388 9436
rect 9688 9380 10416 9408
rect 8792 9296 8876 9324
rect 8988 9296 9072 9352
rect 9156 9324 9240 9380
rect 9324 9352 9380 9380
rect 9660 9352 10444 9380
rect 8512 9240 8596 9296
rect 8820 9268 8876 9296
rect 9016 9268 9072 9296
rect 9184 9296 9240 9324
rect 9352 9296 9380 9352
rect 9632 9324 9940 9352
rect 9632 9296 9688 9324
rect 8820 9240 8904 9268
rect 6524 9184 7000 9212
rect 4340 9156 4872 9184
rect 4928 9156 5124 9184
rect 4340 9128 4956 9156
rect 5012 9128 5124 9156
rect 5404 9128 5460 9184
rect 5600 9156 5740 9184
rect 5628 9128 5684 9156
rect 6020 9128 6412 9184
rect 6496 9156 6944 9184
rect 7280 9156 7476 9212
rect 6468 9128 6888 9156
rect 3864 8568 4228 9128
rect 4340 9100 4648 9128
rect 4788 9100 5124 9128
rect 5376 9100 5460 9128
rect 5600 9100 5656 9128
rect 5992 9100 6860 9128
rect 4340 9072 4564 9100
rect 4872 9072 5096 9100
rect 4312 9016 4508 9072
rect 4984 9044 5096 9072
rect 5012 9016 5096 9044
rect 5348 9072 5516 9100
rect 5600 9072 5628 9100
rect 5964 9072 6356 9100
rect 6412 9072 6860 9100
rect 7308 9072 7476 9156
rect 7560 9128 8008 9240
rect 8540 9184 8624 9240
rect 8848 9184 8904 9240
rect 9016 9212 9100 9268
rect 9184 9240 9268 9296
rect 9352 9268 9408 9296
rect 9044 9184 9100 9212
rect 9212 9212 9268 9240
rect 9380 9212 9408 9268
rect 9604 9268 9688 9296
rect 9744 9296 9884 9324
rect 9744 9268 9856 9296
rect 9604 9240 9828 9268
rect 9576 9212 9800 9240
rect 8568 9128 8652 9184
rect 8876 9128 8932 9184
rect 9044 9128 9128 9184
rect 9212 9156 9296 9212
rect 5348 9016 5600 9072
rect 5964 9044 6888 9072
rect 5936 9016 6888 9044
rect 7308 9016 7504 9072
rect 4312 8680 4480 9016
rect 5012 8680 5068 9016
rect 5348 8988 5572 9016
rect 5320 8904 5376 8988
rect 5460 8960 5572 8988
rect 5908 8960 6888 9016
rect 5320 8848 5348 8904
rect 5516 8848 5544 8960
rect 5880 8932 6888 8960
rect 5852 8904 6888 8932
rect 5852 8876 6244 8904
rect 6272 8876 6888 8904
rect 5320 8736 5544 8848
rect 5824 8848 6216 8876
rect 5824 8820 6188 8848
rect 5796 8792 6188 8820
rect 5768 8764 6160 8792
rect 6272 8764 6300 8876
rect 6356 8848 6888 8876
rect 6384 8792 6888 8848
rect 6412 8764 6888 8792
rect 5768 8736 6132 8764
rect 5320 8708 5376 8736
rect 5348 8680 5376 8708
rect 5544 8680 5572 8736
rect 5740 8708 6132 8736
rect 6244 8736 6384 8764
rect 6440 8736 6888 8764
rect 6244 8708 6888 8736
rect 4312 8624 4508 8680
rect 5012 8652 5096 8680
rect 3864 8540 4256 8568
rect 3892 8428 4256 8540
rect 4340 8540 4508 8624
rect 5040 8596 5096 8652
rect 5348 8624 5404 8680
rect 5572 8652 5600 8680
rect 5712 8652 6104 8708
rect 6244 8680 6468 8708
rect 6496 8680 6888 8708
rect 7336 8680 7504 9016
rect 6216 8652 6468 8680
rect 6552 8652 6888 8680
rect 5516 8624 5600 8652
rect 5684 8624 6076 8652
rect 6216 8624 6244 8652
rect 6328 8624 6468 8652
rect 6608 8624 6860 8652
rect 7308 8624 7504 8680
rect 5376 8596 5404 8624
rect 5488 8596 5628 8624
rect 5040 8540 5124 8596
rect 5376 8568 5432 8596
rect 5460 8568 5656 8596
rect 5684 8568 6048 8624
rect 6188 8596 6216 8624
rect 6160 8568 6216 8596
rect 6384 8568 6440 8624
rect 6720 8596 6804 8624
rect 4340 8484 4536 8540
rect 5068 8512 5124 8540
rect 5404 8540 5628 8568
rect 5656 8540 6020 8568
rect 6104 8540 6244 8568
rect 5404 8512 5600 8540
rect 5684 8512 5992 8540
rect 6076 8512 6272 8540
rect 6356 8512 6412 8568
rect 6692 8540 6776 8596
rect 7308 8540 7476 8624
rect 7588 8568 7952 9128
rect 7980 9100 8008 9128
rect 8596 9100 8652 9128
rect 8596 9072 8680 9100
rect 8904 9072 8960 9128
rect 9072 9100 9128 9128
rect 9240 9128 9296 9156
rect 9408 9156 9436 9212
rect 9576 9184 9856 9212
rect 9576 9156 9912 9184
rect 9408 9128 9464 9156
rect 9576 9128 9772 9156
rect 9828 9128 9940 9156
rect 10024 9128 10080 9352
rect 10164 9324 10444 9352
rect 10220 9296 10360 9324
rect 10388 9296 10472 9324
rect 10248 9268 10360 9296
rect 10416 9268 10472 9296
rect 10276 9240 10500 9268
rect 10248 9212 10500 9240
rect 10220 9184 10528 9212
rect 10164 9156 10304 9184
rect 10136 9128 10248 9156
rect 9240 9100 9324 9128
rect 9072 9072 9156 9100
rect 8624 9044 8680 9072
rect 8932 9044 8988 9072
rect 9100 9044 9156 9072
rect 9268 9072 9324 9100
rect 9436 9072 9464 9128
rect 9268 9044 9352 9072
rect 8624 9016 8708 9044
rect 8932 9016 9016 9044
rect 8652 8988 8708 9016
rect 8960 8988 9016 9016
rect 9100 8988 9184 9044
rect 9296 9016 9352 9044
rect 9464 9016 9492 9072
rect 9548 9016 9744 9128
rect 9884 9100 9996 9128
rect 10024 9100 10220 9128
rect 9912 9072 10164 9100
rect 9968 9016 10136 9072
rect 8652 8960 8736 8988
rect 8960 8960 9044 8988
rect 8680 8932 8736 8960
rect 8988 8932 9044 8960
rect 9128 8932 9212 8988
rect 9296 8960 9380 9016
rect 9492 8988 9520 9016
rect 9548 8988 9772 9016
rect 9912 8988 10192 9016
rect 9492 8960 9548 8988
rect 9324 8932 9408 8960
rect 9520 8932 9548 8960
rect 9576 8932 9772 8988
rect 9884 8960 9996 8988
rect 9828 8932 9968 8960
rect 8680 8904 8764 8932
rect 8988 8904 9072 8932
rect 8708 8876 8792 8904
rect 9016 8876 9072 8904
rect 9156 8904 9212 8932
rect 9352 8904 9408 8932
rect 9548 8904 9912 8932
rect 9156 8876 9240 8904
rect 9352 8876 9436 8904
rect 9548 8876 9884 8904
rect 8736 8848 8792 8876
rect 9044 8848 9100 8876
rect 8736 8820 8820 8848
rect 9044 8820 9128 8848
rect 9184 8820 9268 8876
rect 9380 8848 9436 8876
rect 9576 8848 9716 8876
rect 9744 8848 9828 8876
rect 9380 8820 9464 8848
rect 9604 8820 9688 8848
rect 9744 8820 9856 8848
rect 8764 8792 8820 8820
rect 9072 8792 9128 8820
rect 8764 8764 8848 8792
rect 9072 8764 9156 8792
rect 9212 8764 9296 8820
rect 9408 8792 9492 8820
rect 9604 8792 9912 8820
rect 9436 8764 9520 8792
rect 9632 8764 9996 8792
rect 10024 8764 10080 8988
rect 10108 8960 10220 8988
rect 10332 8960 10528 9184
rect 11144 9156 11200 9716
rect 11228 9688 11284 9716
rect 11704 9688 12068 9716
rect 12152 9688 12656 9744
rect 13328 9716 13384 9744
rect 13776 9716 13832 9744
rect 11228 9660 11312 9688
rect 11732 9660 12040 9688
rect 12124 9660 12488 9688
rect 12572 9660 12656 9688
rect 11228 9632 11424 9660
rect 11760 9632 11984 9660
rect 12124 9632 12460 9660
rect 12628 9632 12712 9660
rect 13300 9632 13328 9716
rect 13692 9688 13776 9716
rect 13888 9688 13916 9772
rect 13356 9660 13664 9688
rect 13888 9660 14224 9688
rect 13860 9632 14420 9660
rect 11228 9604 11508 9632
rect 11228 9576 11592 9604
rect 11228 9548 11648 9576
rect 11788 9548 11956 9632
rect 12096 9604 12460 9632
rect 12488 9604 12572 9632
rect 12712 9604 12768 9632
rect 13244 9604 13328 9632
rect 13804 9604 13916 9632
rect 14140 9604 14560 9632
rect 12096 9576 12432 9604
rect 12488 9576 12656 9604
rect 12768 9576 12796 9604
rect 13160 9576 13328 9604
rect 13748 9576 13916 9604
rect 14364 9576 14672 9604
rect 12068 9548 12432 9576
rect 11228 9520 11676 9548
rect 11228 9492 11704 9520
rect 11760 9492 11984 9548
rect 12068 9520 12404 9548
rect 12460 9520 12740 9576
rect 13104 9548 13440 9576
rect 13608 9548 13944 9576
rect 14504 9548 14784 9576
rect 13048 9520 13216 9548
rect 13244 9520 14224 9548
rect 14616 9520 14868 9548
rect 12040 9492 12404 9520
rect 12432 9492 12740 9520
rect 12992 9492 13132 9520
rect 13244 9492 14420 9520
rect 14728 9492 14952 9520
rect 11228 9464 11928 9492
rect 12040 9464 12376 9492
rect 12432 9464 12712 9492
rect 12936 9464 13076 9492
rect 13244 9464 14560 9492
rect 14812 9464 15008 9492
rect 11228 9436 11788 9464
rect 11984 9436 12376 9464
rect 12404 9436 12712 9464
rect 12908 9436 13020 9464
rect 13244 9436 13972 9464
rect 14308 9436 14672 9464
rect 14896 9436 15092 9464
rect 11228 9408 11648 9436
rect 11844 9408 12348 9436
rect 12404 9408 12684 9436
rect 12852 9408 12964 9436
rect 13188 9408 14000 9436
rect 14476 9408 14784 9436
rect 14952 9408 15148 9436
rect 11228 9380 11508 9408
rect 11704 9380 12348 9408
rect 12376 9380 12684 9408
rect 12824 9380 12936 9408
rect 13132 9380 14000 9408
rect 14588 9380 14868 9408
rect 15036 9380 15204 9408
rect 11228 9352 11396 9380
rect 11564 9352 12320 9380
rect 12376 9352 12656 9380
rect 12796 9352 12908 9380
rect 13048 9352 13216 9380
rect 13272 9352 14000 9380
rect 14700 9352 14924 9380
rect 15092 9352 15260 9380
rect 11228 9324 11340 9352
rect 11424 9324 12320 9352
rect 12348 9324 12600 9352
rect 12768 9324 12880 9352
rect 12992 9324 13132 9352
rect 11228 9156 11312 9324
rect 11368 9296 11816 9324
rect 11340 9184 11396 9296
rect 11480 9268 11676 9296
rect 11928 9268 12292 9324
rect 12348 9296 12460 9324
rect 11480 9240 11564 9268
rect 11732 9240 11900 9268
rect 11928 9240 12264 9268
rect 12320 9240 12460 9296
rect 12740 9296 12852 9324
rect 12964 9296 13048 9324
rect 12740 9268 12824 9296
rect 12908 9268 12992 9296
rect 13300 9268 14028 9352
rect 14812 9324 15008 9352
rect 15148 9324 15288 9352
rect 14896 9296 15064 9324
rect 15204 9296 15344 9324
rect 14980 9268 15148 9296
rect 15260 9268 15372 9296
rect 12712 9240 12796 9268
rect 12880 9240 12936 9268
rect 13328 9240 14028 9268
rect 15036 9240 15148 9268
rect 15288 9240 15428 9268
rect 11480 9212 11536 9240
rect 11592 9212 12264 9240
rect 12292 9212 12460 9240
rect 12516 9212 12768 9240
rect 11480 9184 11508 9212
rect 11564 9184 12236 9212
rect 12292 9184 12768 9212
rect 13328 9184 14056 9240
rect 15344 9212 15456 9240
rect 15372 9184 15512 9212
rect 11368 9156 11508 9184
rect 11144 9100 11172 9156
rect 10164 8932 10276 8960
rect 10304 8932 10528 8960
rect 10192 8904 10500 8932
rect 10248 8848 10500 8904
rect 10220 8820 10472 8848
rect 10192 8792 10332 8820
rect 10388 8792 10472 8820
rect 11116 8792 11172 9100
rect 11228 9100 11340 9156
rect 11396 9100 11508 9156
rect 11536 9156 12236 9184
rect 11536 9128 12208 9156
rect 12264 9128 12740 9184
rect 11564 9100 12208 9128
rect 12236 9100 12740 9128
rect 13356 9156 14056 9184
rect 15428 9156 15540 9184
rect 13356 9128 14084 9156
rect 15456 9128 15568 9156
rect 13356 9100 13552 9128
rect 13944 9100 14084 9128
rect 15484 9100 15596 9128
rect 11228 9072 11368 9100
rect 11424 9072 11536 9100
rect 11228 9044 11396 9072
rect 11452 9044 11536 9072
rect 11592 9044 12180 9100
rect 12208 9044 12712 9100
rect 13356 9072 13524 9100
rect 13972 9072 14084 9100
rect 15512 9072 15624 9100
rect 11228 9016 11424 9044
rect 11480 9016 11564 9044
rect 11620 9016 12152 9044
rect 11228 8932 11312 9016
rect 11340 8988 11452 9016
rect 11508 8988 11592 9016
rect 11648 8988 12152 9016
rect 12180 9016 12712 9044
rect 12180 8988 12404 9016
rect 11340 8960 11480 8988
rect 11200 8904 11312 8932
rect 11368 8932 11480 8960
rect 11536 8960 11620 8988
rect 11536 8932 11648 8960
rect 11676 8932 12124 8988
rect 12152 8932 12376 8988
rect 11368 8904 11508 8932
rect 11564 8904 11648 8932
rect 11704 8904 12096 8932
rect 11200 8792 11340 8904
rect 10108 8764 10444 8792
rect 11144 8764 11340 8792
rect 8792 8736 8848 8764
rect 9100 8736 9156 8764
rect 9240 8736 9324 8764
rect 9436 8736 9548 8764
rect 9660 8736 10416 8764
rect 11172 8736 11340 8764
rect 8792 8708 8876 8736
rect 8820 8680 8876 8708
rect 9128 8708 9184 8736
rect 9268 8708 9352 8736
rect 9464 8708 9576 8736
rect 9688 8708 10388 8736
rect 9128 8680 9212 8708
rect 8820 8652 8904 8680
rect 9156 8652 9212 8680
rect 9296 8680 9352 8708
rect 9492 8680 9604 8708
rect 9716 8680 10360 8708
rect 11228 8680 11340 8736
rect 11368 8876 11536 8904
rect 11592 8876 11676 8904
rect 11732 8876 12096 8904
rect 12124 8876 12348 8932
rect 12572 8904 12712 9016
rect 13384 9044 13524 9072
rect 13580 9044 13916 9072
rect 13972 9044 14112 9072
rect 15540 9044 15652 9072
rect 13384 8988 13552 9044
rect 13580 9016 13888 9044
rect 13608 8988 13888 9016
rect 13944 8988 14112 9044
rect 15568 9016 15680 9044
rect 15596 8988 15708 9016
rect 13412 8932 13580 8988
rect 13608 8960 13860 8988
rect 13916 8960 14140 8988
rect 15624 8960 15736 8988
rect 13636 8932 13860 8960
rect 13412 8904 13608 8932
rect 11368 8848 11564 8876
rect 11620 8848 12068 8876
rect 11368 8820 11592 8848
rect 11648 8820 12068 8848
rect 12096 8848 12320 8876
rect 12096 8820 12292 8848
rect 11368 8764 11620 8820
rect 11676 8764 12040 8820
rect 12068 8792 12292 8820
rect 12600 8792 12712 8904
rect 13440 8848 13636 8904
rect 13664 8876 13832 8932
rect 13888 8904 14140 8960
rect 15652 8932 15764 8960
rect 15680 8904 15792 8932
rect 13692 8848 13804 8876
rect 13860 8848 14168 8904
rect 15708 8876 15792 8904
rect 15736 8848 15820 8876
rect 13440 8792 13664 8848
rect 13692 8820 13776 8848
rect 13832 8820 14168 8848
rect 13720 8792 13776 8820
rect 13804 8792 14168 8820
rect 15764 8820 15848 8848
rect 15764 8792 15876 8820
rect 12068 8764 12264 8792
rect 11368 8736 12012 8764
rect 11368 8708 11620 8736
rect 11648 8708 12012 8736
rect 12040 8708 12264 8764
rect 12628 8764 12712 8792
rect 12628 8708 12740 8764
rect 13468 8736 13692 8792
rect 13804 8764 14196 8792
rect 15792 8764 15876 8792
rect 13776 8736 14196 8764
rect 13468 8708 14196 8736
rect 15820 8708 15904 8764
rect 11368 8680 11564 8708
rect 9296 8652 9380 8680
rect 9520 8652 9632 8680
rect 9772 8652 10332 8680
rect 11256 8652 11312 8680
rect 11340 8652 11508 8680
rect 11620 8652 11984 8708
rect 12012 8680 12292 8708
rect 12012 8652 12348 8680
rect 12656 8652 12740 8708
rect 8848 8624 8932 8652
rect 9156 8624 9240 8652
rect 9324 8624 9408 8652
rect 9576 8624 9660 8652
rect 9800 8624 10276 8652
rect 11256 8624 11452 8652
rect 8876 8596 8932 8624
rect 9184 8596 9240 8624
rect 9352 8596 9436 8624
rect 9604 8596 9716 8624
rect 9884 8596 10220 8624
rect 11592 8596 11956 8652
rect 11984 8624 12404 8652
rect 11984 8596 12432 8624
rect 12656 8596 12768 8652
rect 13496 8624 14224 8708
rect 15848 8652 15932 8708
rect 8876 8568 8960 8596
rect 6692 8512 6748 8540
rect 5068 8484 5152 8512
rect 5432 8484 5544 8512
rect 5712 8484 5992 8512
rect 6020 8484 6076 8512
rect 6132 8484 6272 8512
rect 6328 8484 6384 8512
rect 6664 8484 6748 8512
rect 7280 8484 7476 8540
rect 7560 8540 7952 8568
rect 8904 8540 8960 8568
rect 9212 8568 9268 8596
rect 9380 8568 9464 8596
rect 9660 8568 9772 8596
rect 9996 8568 10108 8596
rect 11564 8568 11928 8596
rect 11956 8568 12488 8596
rect 12684 8568 12768 8596
rect 9212 8540 9296 8568
rect 9408 8540 9520 8568
rect 9688 8540 9828 8568
rect 11564 8540 11900 8568
rect 11956 8540 12544 8568
rect 4368 8428 4536 8484
rect 5096 8456 5152 8484
rect 5460 8456 5516 8484
rect 5096 8428 5180 8456
rect 5488 8428 5544 8456
rect 5684 8428 6020 8484
rect 6132 8456 6356 8484
rect 6664 8456 6720 8484
rect 6160 8428 6328 8456
rect 6636 8428 6720 8456
rect 7280 8428 7448 8484
rect 7560 8428 7924 8540
rect 8904 8512 8988 8540
rect 9240 8512 9296 8540
rect 9436 8512 9548 8540
rect 9744 8512 9912 8540
rect 11536 8512 11900 8540
rect 11928 8512 12600 8540
rect 12684 8512 12796 8568
rect 13524 8540 14252 8624
rect 15876 8596 15960 8652
rect 15904 8540 15988 8596
rect 13524 8512 14280 8540
rect 8932 8484 8988 8512
rect 9268 8484 9324 8512
rect 9464 8484 9604 8512
rect 9828 8484 10024 8512
rect 11536 8484 11872 8512
rect 11928 8484 12152 8512
rect 12208 8484 12628 8512
rect 12684 8484 12824 8512
rect 8960 8456 9016 8484
rect 9268 8456 9352 8484
rect 9520 8456 9632 8484
rect 9912 8456 10108 8484
rect 8960 8428 9044 8456
rect 9296 8428 9352 8456
rect 9548 8428 9716 8456
rect 10052 8428 10108 8456
rect 11508 8456 11872 8484
rect 11508 8428 11844 8456
rect 11900 8428 12124 8484
rect 12264 8456 12824 8484
rect 12292 8428 12852 8456
rect 13552 8428 14280 8512
rect 3892 8400 4284 8428
rect 3920 8344 4284 8400
rect 4368 8372 4564 8428
rect 5124 8400 5180 8428
rect 5516 8400 5572 8428
rect 5124 8372 5208 8400
rect 5544 8372 5628 8400
rect 5656 8372 5796 8428
rect 4396 8344 4564 8372
rect 5152 8344 5236 8372
rect 5572 8344 5768 8372
rect 5908 8344 6048 8428
rect 6188 8400 6300 8428
rect 6636 8400 6692 8428
rect 6188 8372 6272 8400
rect 6608 8372 6692 8400
rect 7252 8372 7448 8428
rect 7532 8400 7924 8428
rect 8988 8400 9044 8428
rect 6160 8344 6244 8372
rect 6580 8344 6664 8372
rect 7252 8344 7420 8372
rect 7532 8344 7896 8400
rect 8988 8372 9072 8400
rect 9324 8372 9380 8428
rect 9604 8400 9772 8428
rect 11480 8400 11844 8428
rect 9660 8372 9856 8400
rect 11480 8372 11816 8400
rect 11872 8372 12096 8428
rect 12348 8400 12880 8428
rect 12404 8372 12908 8400
rect 9016 8344 9072 8372
rect 9352 8344 9408 8372
rect 9744 8344 9968 8372
rect 11452 8344 11816 8372
rect 11844 8344 12096 8372
rect 12460 8344 12964 8372
rect 13580 8344 14308 8428
rect 3920 8288 4312 8344
rect 4396 8288 4592 8344
rect 5180 8316 5236 8344
rect 5628 8316 5768 8344
rect 5936 8316 6048 8344
rect 6076 8316 6188 8344
rect 6580 8316 6636 8344
rect 5180 8288 5264 8316
rect 5684 8288 5880 8316
rect 5908 8288 6132 8316
rect 6552 8288 6636 8316
rect 7224 8288 7420 8344
rect 7504 8288 7896 8344
rect 9044 8316 9100 8344
rect 9044 8288 9128 8316
rect 9380 8288 9436 8344
rect 9828 8316 10052 8344
rect 9940 8288 10052 8316
rect 11424 8288 11788 8344
rect 11844 8316 12068 8344
rect 12516 8316 12992 8344
rect 11816 8288 12068 8316
rect 12544 8288 13048 8316
rect 3948 8260 4312 8288
rect 3948 8176 4340 8260
rect 4424 8232 4620 8288
rect 5208 8260 5292 8288
rect 5796 8260 6020 8288
rect 6524 8260 6608 8288
rect 5236 8232 5320 8260
rect 6496 8232 6580 8260
rect 7196 8232 7392 8288
rect 7504 8260 7868 8288
rect 9072 8260 9128 8288
rect 9408 8260 9464 8288
rect 4424 8204 4648 8232
rect 5264 8204 5348 8232
rect 6468 8204 6552 8232
rect 4452 8176 4648 8204
rect 5292 8176 5376 8204
rect 6440 8176 6580 8204
rect 7168 8176 7364 8232
rect 7476 8204 7868 8260
rect 9100 8232 9156 8260
rect 9100 8204 9184 8232
rect 9436 8204 9492 8260
rect 11396 8232 11760 8288
rect 11816 8260 12040 8288
rect 12544 8260 13104 8288
rect 13608 8260 14336 8344
rect 3976 8120 4368 8176
rect 4452 8148 4676 8176
rect 4480 8120 4676 8148
rect 5320 8148 5432 8176
rect 6384 8148 6608 8176
rect 7140 8148 7364 8176
rect 7448 8176 7868 8204
rect 9128 8176 9184 8204
rect 9464 8176 9520 8204
rect 11368 8176 11732 8232
rect 11788 8204 12040 8260
rect 12516 8232 13188 8260
rect 13608 8232 14364 8260
rect 12516 8204 13272 8232
rect 5320 8120 5460 8148
rect 6356 8120 6496 8148
rect 6524 8120 6636 8148
rect 7140 8120 7336 8148
rect 7448 8120 7840 8176
rect 9156 8148 9212 8176
rect 9156 8120 9240 8148
rect 11340 8120 11704 8176
rect 11760 8148 12012 8204
rect 12516 8148 12628 8204
rect 11732 8120 12012 8148
rect 4004 8064 4396 8120
rect 4480 8092 4704 8120
rect 5320 8092 5516 8120
rect 6300 8092 6412 8120
rect 6440 8092 6524 8120
rect 6552 8092 6636 8120
rect 7112 8092 7336 8120
rect 4508 8064 4704 8092
rect 5292 8064 5376 8092
rect 5404 8064 5572 8092
rect 6244 8064 6384 8092
rect 6468 8064 6552 8092
rect 6580 8064 6664 8092
rect 7112 8064 7308 8092
rect 7420 8064 7812 8120
rect 9184 8092 9240 8120
rect 4004 8036 4424 8064
rect 4508 8036 4732 8064
rect 5264 8036 5348 8064
rect 5376 8036 5460 8064
rect 5488 8036 5656 8064
rect 6160 8036 6328 8064
rect 6468 8036 6692 8064
rect 7084 8036 7308 8064
rect 7392 8036 7812 8064
rect 9212 8036 9268 8092
rect 11312 8064 11676 8120
rect 11732 8092 11984 8120
rect 4032 8008 4424 8036
rect 4536 8008 4760 8036
rect 5264 8008 5460 8036
rect 5544 8008 5768 8036
rect 6048 8008 6272 8036
rect 6496 8008 6580 8036
rect 6608 8008 6720 8036
rect 7056 8008 7280 8036
rect 7392 8008 7784 8036
rect 9240 8008 9296 8036
rect 11284 8008 11648 8064
rect 11704 8036 11984 8092
rect 12488 8064 12628 8148
rect 12684 8176 13440 8204
rect 13636 8176 14364 8232
rect 15652 8176 15848 8204
rect 12684 8148 14392 8176
rect 15092 8148 15848 8176
rect 12684 8120 15820 8148
rect 12684 8092 15344 8120
rect 12712 8064 12908 8092
rect 12964 8064 14588 8092
rect 4032 7980 4452 8008
rect 4060 7924 4480 7980
rect 4564 7952 4788 8008
rect 5236 7980 5320 8008
rect 5348 7980 5432 8008
rect 5628 7980 6188 8008
rect 6524 7980 6608 8008
rect 6636 7980 6748 8008
rect 5208 7952 5292 7980
rect 5320 7952 5404 7980
rect 5712 7952 6104 7980
rect 6552 7952 6636 7980
rect 6664 7952 6776 7980
rect 7028 7952 7252 8008
rect 7364 7980 7784 8008
rect 4592 7924 4816 7952
rect 5180 7924 5404 7952
rect 6552 7924 6804 7952
rect 7000 7924 7224 7952
rect 7336 7924 7756 7980
rect 9268 7952 9324 8008
rect 11256 7952 11620 8008
rect 11676 7980 11956 8036
rect 11648 7952 11956 7980
rect 12488 7952 12656 8064
rect 12712 7980 12936 8064
rect 13020 8036 14644 8064
rect 13076 8008 14784 8036
rect 13132 7980 14812 8008
rect 12740 7952 12936 7980
rect 13160 7952 14868 7980
rect 4088 7896 4508 7924
rect 4620 7896 4844 7924
rect 5180 7896 5264 7924
rect 5292 7896 5376 7924
rect 6580 7896 6664 7924
rect 6692 7896 6916 7924
rect 6972 7896 7196 7924
rect 7308 7896 7728 7924
rect 11228 7896 11592 7952
rect 11648 7924 11928 7952
rect 4088 7868 4536 7896
rect 4620 7868 4872 7896
rect 5124 7868 5236 7896
rect 5264 7868 5348 7896
rect 4116 7840 4536 7868
rect 4648 7840 4900 7868
rect 5068 7840 5348 7868
rect 6608 7868 6692 7896
rect 6720 7868 7196 7896
rect 7280 7868 7728 7896
rect 4116 7812 4564 7840
rect 4676 7812 5208 7840
rect 5236 7812 5320 7840
rect 6608 7812 6720 7868
rect 6748 7840 7168 7868
rect 7280 7840 7700 7868
rect 11200 7840 11564 7896
rect 11620 7868 11928 7924
rect 12516 7868 12684 7952
rect 12740 7868 12964 7952
rect 13216 7924 14896 7952
rect 13272 7896 14924 7924
rect 13272 7868 14952 7896
rect 11620 7840 11844 7868
rect 12516 7840 12712 7868
rect 6748 7812 7140 7840
rect 7252 7812 7700 7840
rect 4144 7784 4592 7812
rect 4704 7784 5180 7812
rect 5208 7784 5320 7812
rect 6636 7784 6748 7812
rect 6776 7784 7112 7812
rect 7224 7784 7672 7812
rect 11172 7784 11536 7840
rect 11592 7812 11732 7840
rect 11564 7784 11648 7812
rect 4172 7756 4620 7784
rect 4732 7756 5152 7784
rect 4172 7728 4648 7756
rect 4760 7728 5152 7756
rect 5180 7728 5292 7784
rect 6636 7756 7084 7784
rect 7196 7756 7644 7784
rect 4200 7700 4648 7728
rect 4788 7700 5124 7728
rect 5152 7700 5292 7728
rect 4200 7672 4676 7700
rect 4816 7672 5292 7700
rect 4228 7644 4704 7672
rect 4844 7644 5292 7672
rect 4256 7616 4732 7644
rect 4872 7616 5292 7644
rect 6608 7728 7056 7756
rect 7168 7728 7644 7756
rect 11144 7728 11508 7784
rect 12544 7756 12712 7840
rect 12768 7840 12964 7868
rect 13300 7840 14952 7868
rect 12768 7756 12992 7840
rect 13300 7812 14980 7840
rect 13328 7784 15008 7812
rect 13328 7756 16072 7784
rect 12544 7728 12740 7756
rect 6608 7700 7028 7728
rect 7168 7700 7616 7728
rect 6608 7672 7000 7700
rect 7140 7672 7616 7700
rect 11116 7672 11480 7728
rect 6608 7644 6972 7672
rect 7112 7644 7588 7672
rect 6608 7616 6944 7644
rect 7084 7616 7560 7644
rect 11088 7616 11452 7672
rect 12572 7644 12740 7728
rect 12796 7728 12992 7756
rect 13356 7728 16072 7756
rect 12796 7672 13020 7728
rect 13356 7700 14924 7728
rect 12824 7644 13020 7672
rect 13384 7672 14924 7700
rect 13384 7644 14896 7672
rect 4284 7588 4760 7616
rect 4900 7588 5292 7616
rect 6580 7588 6916 7616
rect 7056 7588 7532 7616
rect 11060 7588 11424 7616
rect 4284 7560 4816 7588
rect 4928 7560 5320 7588
rect 6524 7560 6888 7588
rect 7000 7560 7532 7588
rect 11032 7560 11424 7588
rect 12600 7560 12768 7644
rect 12824 7560 13048 7644
rect 13412 7616 13776 7644
rect 13244 7588 13580 7616
rect 13748 7588 13776 7616
rect 13860 7588 14868 7644
rect 13160 7560 13300 7588
rect 13496 7560 13552 7588
rect 13748 7560 13804 7588
rect 4312 7532 4844 7560
rect 4984 7532 5348 7560
rect 6468 7532 6832 7560
rect 6972 7532 7504 7560
rect 11032 7532 11396 7560
rect 12600 7532 12796 7560
rect 4340 7504 4872 7532
rect 5012 7504 5404 7532
rect 6412 7504 6804 7532
rect 6944 7504 7476 7532
rect 11004 7504 11396 7532
rect 4368 7476 4900 7504
rect 5068 7476 5488 7504
rect 6328 7476 6748 7504
rect 6916 7476 7448 7504
rect 11004 7476 11368 7504
rect 4396 7448 4956 7476
rect 5124 7448 5600 7476
rect 6216 7448 6692 7476
rect 6860 7448 7420 7476
rect 9828 7448 10080 7476
rect 10976 7448 11368 7476
rect 12628 7448 12796 7532
rect 12852 7532 13048 7560
rect 13076 7532 13188 7560
rect 12852 7504 13132 7532
rect 12852 7476 13076 7504
rect 13524 7476 13580 7560
rect 12852 7448 13048 7476
rect 13552 7448 13580 7476
rect 4424 7420 4984 7448
rect 5152 7420 5768 7448
rect 6048 7420 6664 7448
rect 6832 7420 7392 7448
rect 9576 7420 10332 7448
rect 10976 7420 11340 7448
rect 12628 7420 12824 7448
rect 4452 7392 5040 7420
rect 5208 7392 6608 7420
rect 6776 7392 7364 7420
rect 9436 7392 9856 7420
rect 10052 7392 10500 7420
rect 10948 7392 11340 7420
rect 4480 7364 5096 7392
rect 5292 7364 6524 7392
rect 6720 7364 7336 7392
rect 9352 7364 9604 7392
rect 10304 7364 10612 7392
rect 10948 7364 11312 7392
rect 4508 7336 5124 7364
rect 5348 7336 6468 7364
rect 6692 7336 7308 7364
rect 9268 7336 9492 7364
rect 10444 7336 10696 7364
rect 10920 7336 11312 7364
rect 4536 7308 5180 7336
rect 5432 7308 6384 7336
rect 6636 7308 7280 7336
rect 9184 7308 9380 7336
rect 10556 7308 10780 7336
rect 10920 7308 11284 7336
rect 12656 7308 12824 7420
rect 12880 7420 13020 7448
rect 12880 7392 12992 7420
rect 13524 7392 13580 7448
rect 13776 7392 13804 7560
rect 13860 7560 15988 7588
rect 13860 7532 15960 7560
rect 13832 7476 14924 7504
rect 12880 7364 12964 7392
rect 13524 7364 13552 7392
rect 12880 7308 12936 7364
rect 13412 7336 13552 7364
rect 13748 7336 13804 7392
rect 14812 7364 14868 7392
rect 13832 7336 15988 7364
rect 13300 7308 13776 7336
rect 4564 7280 5264 7308
rect 5544 7280 6272 7308
rect 6552 7280 7252 7308
rect 9128 7280 9296 7308
rect 10668 7280 10864 7308
rect 10892 7280 11256 7308
rect 4592 7252 5320 7280
rect 5712 7252 6104 7280
rect 6496 7252 7224 7280
rect 9072 7252 9212 7280
rect 10752 7252 11256 7280
rect 4620 7224 5404 7252
rect 6412 7224 7196 7252
rect 9044 7224 9156 7252
rect 10836 7224 11228 7252
rect 4676 7196 5516 7224
rect 6300 7196 7140 7224
rect 9044 7196 9128 7224
rect 10864 7196 11228 7224
rect 12684 7224 12796 7308
rect 12880 7280 12908 7308
rect 13244 7280 13412 7308
rect 13664 7280 13776 7308
rect 14812 7308 15988 7336
rect 12852 7252 12908 7280
rect 13188 7252 13328 7280
rect 13636 7252 13720 7280
rect 14812 7252 14868 7308
rect 12852 7224 12880 7252
rect 13160 7224 13272 7252
rect 13636 7224 13692 7252
rect 14196 7224 14252 7252
rect 14448 7224 14532 7252
rect 12684 7196 12768 7224
rect 4704 7168 5628 7196
rect 6188 7168 7112 7196
rect 9072 7168 9212 7196
rect 4732 7140 7084 7168
rect 9100 7140 9352 7168
rect 10836 7140 11200 7196
rect 4788 7112 7028 7140
rect 9156 7112 9912 7140
rect 10808 7112 11200 7140
rect 12712 7112 12768 7196
rect 4844 7084 6972 7112
rect 9100 7084 10136 7112
rect 10808 7084 11256 7112
rect 12740 7084 12768 7112
rect 12824 7168 12880 7224
rect 13132 7196 13216 7224
rect 13132 7168 13188 7196
rect 13608 7168 13664 7224
rect 13888 7196 13972 7224
rect 14196 7196 14280 7224
rect 14448 7196 14560 7224
rect 4872 7056 6944 7084
rect 9044 7056 10304 7084
rect 10780 7056 11284 7084
rect 4928 7028 6888 7056
rect 8988 7028 10416 7056
rect 10780 7028 11144 7056
rect 11200 7028 11312 7056
rect 12740 7028 12768 7056
rect 4984 7000 6832 7028
rect 8932 7000 10528 7028
rect 5040 6972 6776 7000
rect 8876 6972 10612 7000
rect 10752 6972 11116 7028
rect 11256 7000 11368 7028
rect 11284 6972 11396 7000
rect 5096 6944 6720 6972
rect 8820 6944 10696 6972
rect 10724 6944 11088 6972
rect 11340 6944 11424 6972
rect 5180 6916 6636 6944
rect 8792 6916 11088 6944
rect 11368 6916 11452 6944
rect 12824 6916 12852 7168
rect 13104 7140 13188 7168
rect 13104 7084 13160 7140
rect 13104 6972 13188 7084
rect 13580 6972 13636 7168
rect 13888 7140 14000 7196
rect 14196 7168 14308 7196
rect 14448 7168 14588 7196
rect 14196 7140 14336 7168
rect 14476 7140 14616 7168
rect 13916 7112 14028 7140
rect 14224 7112 14336 7140
rect 14504 7112 14616 7140
rect 14840 7112 14896 7252
rect 13916 7084 14056 7112
rect 13944 7056 14056 7084
rect 14252 7056 14364 7112
rect 14532 7056 14616 7112
rect 14868 7056 14924 7112
rect 13972 7028 14056 7056
rect 14308 7028 14336 7056
rect 14868 7028 15008 7056
rect 14028 7000 14056 7028
rect 14868 7000 16044 7028
rect 14672 6972 15288 7000
rect 13104 6944 13216 6972
rect 5264 6888 6552 6916
rect 8736 6888 11060 6916
rect 11396 6888 11480 6916
rect 5348 6860 6468 6888
rect 8708 6860 9744 6888
rect 10136 6860 11060 6888
rect 11424 6860 11508 6888
rect 12824 6860 12880 6916
rect 13132 6888 13216 6944
rect 13608 6888 13664 6972
rect 14392 6944 14616 6972
rect 14896 6944 14952 6972
rect 14112 6916 14336 6944
rect 14924 6916 14980 6944
rect 13832 6888 14056 6916
rect 14924 6888 15008 6916
rect 5460 6832 6356 6860
rect 8652 6832 9576 6860
rect 10304 6832 11032 6860
rect 11452 6832 11536 6860
rect 12852 6832 12880 6860
rect 13160 6832 13244 6888
rect 13636 6860 13776 6888
rect 14308 6860 14364 6888
rect 14560 6860 14644 6888
rect 14952 6860 15008 6888
rect 13636 6832 13692 6860
rect 5628 6804 6188 6832
rect 8624 6804 9464 6832
rect 10416 6804 11032 6832
rect 11480 6804 11564 6832
rect 12852 6804 12908 6832
rect 13188 6804 13272 6832
rect 13608 6804 13692 6832
rect 8596 6776 9380 6804
rect 10500 6776 11032 6804
rect 11508 6776 11592 6804
rect 12880 6776 12908 6804
rect 13216 6776 13356 6804
rect 13524 6776 13692 6804
rect 8568 6748 9296 6776
rect 9632 6748 10220 6776
rect 10584 6748 11088 6776
rect 11536 6748 11620 6776
rect 12880 6748 12936 6776
rect 13272 6748 13692 6776
rect 14000 6804 14084 6860
rect 14280 6832 14392 6860
rect 14560 6832 14672 6860
rect 14980 6832 15036 6860
rect 14280 6804 14420 6832
rect 14560 6804 14700 6832
rect 14980 6804 15064 6832
rect 14000 6776 14112 6804
rect 14308 6776 14420 6804
rect 14588 6776 14700 6804
rect 15008 6776 15064 6804
rect 14000 6748 14140 6776
rect 8512 6720 9212 6748
rect 9520 6720 10360 6748
rect 10612 6720 11144 6748
rect 11564 6720 11648 6748
rect 12908 6720 12964 6748
rect 13356 6720 13496 6748
rect 8484 6692 9156 6720
rect 9408 6692 10444 6720
rect 10584 6692 11172 6720
rect 8456 6664 9100 6692
rect 9324 6664 10528 6692
rect 10584 6664 11200 6692
rect 11592 6664 11676 6720
rect 12908 6692 12992 6720
rect 13636 6692 13692 6748
rect 14028 6720 14168 6748
rect 14336 6720 14448 6776
rect 14616 6720 14728 6776
rect 15036 6748 15092 6776
rect 15036 6720 15120 6748
rect 14056 6692 14168 6720
rect 14364 6692 14448 6720
rect 14644 6692 14728 6720
rect 15064 6692 15120 6720
rect 12936 6664 13020 6692
rect 13636 6664 13720 6692
rect 14084 6664 14168 6692
rect 14420 6664 14448 6692
rect 15092 6664 15148 6692
rect 8428 6636 9072 6664
rect 9268 6636 11256 6664
rect 11620 6636 11704 6664
rect 12824 6636 12852 6664
rect 12964 6636 13048 6664
rect 8400 6608 9016 6636
rect 9212 6608 11284 6636
rect 11648 6608 11732 6636
rect 8372 6580 8960 6608
rect 9156 6580 9744 6608
rect 8344 6552 8932 6580
rect 9100 6552 9660 6580
rect 9940 6552 9996 6608
rect 10136 6580 11312 6608
rect 11676 6580 11732 6608
rect 12824 6608 12880 6636
rect 13020 6608 13076 6636
rect 13664 6608 13720 6664
rect 15092 6636 15176 6664
rect 15064 6608 15176 6636
rect 12824 6580 12908 6608
rect 13048 6580 13132 6608
rect 13664 6580 13748 6608
rect 14672 6580 15204 6608
rect 1260 6524 2044 6552
rect 2492 6524 2772 6552
rect 2968 6524 3248 6552
rect 3528 6524 3808 6552
rect 4032 6524 4312 6552
rect 4564 6524 4872 6552
rect 8316 6524 8904 6552
rect 9044 6524 9492 6552
rect 1596 6496 2464 6524
rect 1792 6412 2464 6496
rect 1764 6356 2436 6412
rect 2632 6384 2828 6524
rect 2632 6356 2800 6384
rect 3108 6356 3416 6524
rect 3668 6496 3976 6524
rect 3780 6440 3976 6496
rect 3780 6412 3948 6440
rect 1988 6244 2184 6356
rect 2604 6244 2800 6356
rect 1988 6216 2156 6244
rect 2604 6216 2772 6244
rect 3080 6216 3416 6356
rect 3752 6300 3948 6412
rect 4144 6356 4340 6524
rect 4704 6496 4956 6524
rect 8316 6496 8848 6524
rect 9016 6496 9408 6524
rect 4760 6468 4956 6496
rect 8288 6468 8820 6496
rect 8960 6468 9380 6496
rect 4732 6412 4928 6468
rect 8260 6440 8792 6468
rect 8932 6440 9296 6468
rect 9352 6440 9380 6468
rect 8232 6412 8764 6440
rect 8904 6412 9240 6440
rect 4704 6356 4900 6412
rect 8204 6384 8736 6412
rect 8848 6384 9184 6412
rect 9212 6384 9268 6412
rect 9352 6384 9408 6440
rect 8204 6356 8708 6384
rect 8820 6356 9128 6384
rect 9240 6356 9296 6384
rect 4172 6300 4340 6356
rect 4676 6300 4872 6356
rect 8176 6328 8680 6356
rect 8792 6328 9100 6356
rect 9268 6328 9352 6356
rect 9380 6328 9408 6384
rect 8148 6300 8652 6328
rect 8764 6300 9044 6328
rect 9296 6300 9408 6328
rect 3752 6272 3920 6300
rect 1960 6104 2156 6216
rect 2576 6104 2772 6216
rect 3052 6188 3416 6216
rect 3052 6160 3248 6188
rect 3052 6104 3220 6160
rect 1960 6076 2128 6104
rect 1932 5964 2128 6076
rect 2548 5992 2744 6104
rect 3024 5992 3220 6104
rect 2548 5964 2716 5992
rect 3024 5964 3192 5992
rect 1932 5936 2100 5964
rect 1904 5852 2100 5936
rect 2520 5852 2716 5964
rect 2996 5852 3192 5964
rect 3276 5852 3416 6188
rect 3724 6160 3920 6272
rect 3696 6048 3892 6160
rect 3696 6020 3864 6048
rect 3668 5908 3864 6020
rect 4172 5992 4368 6300
rect 4676 6272 4844 6300
rect 8148 6272 8624 6300
rect 8736 6272 9016 6300
rect 9352 6272 9436 6300
rect 4648 6244 4844 6272
rect 8120 6244 8596 6272
rect 8708 6244 9072 6272
rect 9380 6244 9436 6272
rect 4648 6216 4816 6244
rect 4620 6188 4816 6216
rect 8092 6216 8568 6244
rect 8680 6216 8960 6244
rect 9016 6216 9100 6244
rect 9380 6216 9464 6244
rect 8092 6188 8540 6216
rect 8652 6188 8932 6216
rect 9072 6188 9156 6216
rect 9408 6188 9520 6216
rect 4620 6160 4788 6188
rect 4592 6132 4788 6160
rect 8064 6132 8512 6188
rect 8652 6160 8904 6188
rect 9100 6160 9184 6188
rect 8624 6132 8876 6160
rect 9156 6132 9240 6160
rect 9408 6132 9436 6188
rect 9464 6160 9548 6188
rect 9604 6160 9632 6552
rect 9968 6496 9996 6552
rect 10192 6552 10248 6580
rect 10276 6552 10892 6580
rect 10948 6552 11340 6580
rect 11676 6552 11760 6580
rect 12852 6552 12964 6580
rect 13076 6552 13188 6580
rect 13636 6552 13776 6580
rect 14280 6552 15008 6580
rect 10192 6524 10220 6552
rect 10304 6524 10360 6552
rect 10388 6524 10892 6552
rect 10976 6524 11396 6552
rect 11704 6524 11788 6552
rect 9968 6440 10024 6496
rect 10192 6468 10248 6524
rect 10276 6496 10332 6524
rect 10444 6496 10864 6524
rect 11004 6496 11424 6524
rect 11732 6496 11788 6524
rect 12852 6524 12992 6552
rect 13104 6524 13244 6552
rect 13552 6524 13664 6552
rect 13720 6524 13804 6552
rect 13888 6524 14812 6552
rect 12852 6496 13048 6524
rect 13104 6496 13608 6524
rect 13748 6496 14840 6524
rect 10276 6468 10304 6496
rect 10192 6440 10304 6468
rect 10472 6468 10892 6496
rect 11060 6468 11452 6496
rect 11732 6468 11816 6496
rect 10472 6440 10948 6468
rect 11088 6440 11480 6468
rect 11760 6440 11816 6468
rect 9996 6384 10024 6440
rect 10220 6384 10276 6440
rect 10444 6412 10976 6440
rect 11116 6412 11508 6440
rect 11760 6412 11844 6440
rect 10444 6384 11004 6412
rect 11144 6384 11508 6412
rect 11788 6384 11844 6412
rect 12880 6384 13076 6496
rect 13104 6468 13468 6496
rect 13776 6468 14364 6496
rect 14420 6468 14896 6496
rect 13132 6440 13328 6468
rect 13748 6440 13944 6468
rect 13972 6440 14336 6468
rect 14448 6440 14784 6468
rect 14840 6440 14952 6468
rect 9996 6300 10052 6384
rect 10192 6356 10248 6384
rect 10164 6300 10248 6356
rect 10416 6356 11032 6384
rect 11172 6356 11536 6384
rect 11788 6356 11872 6384
rect 10416 6328 11060 6356
rect 11200 6328 11564 6356
rect 11816 6328 11872 6356
rect 10024 6244 10052 6300
rect 10136 6272 10192 6300
rect 10024 6216 10080 6244
rect 10108 6216 10164 6272
rect 10024 6188 10136 6216
rect 10220 6188 10276 6300
rect 10388 6272 10780 6328
rect 10808 6300 11088 6328
rect 11228 6300 11592 6328
rect 11816 6300 11900 6328
rect 12908 6300 13104 6384
rect 13132 6356 13356 6440
rect 13720 6384 13916 6440
rect 14000 6412 14364 6440
rect 14420 6412 14756 6440
rect 14840 6412 14980 6440
rect 14000 6384 14784 6412
rect 14840 6384 15008 6412
rect 13692 6356 13944 6384
rect 13972 6356 15036 6384
rect 10836 6272 11116 6300
rect 11256 6272 11620 6300
rect 10360 6244 10752 6272
rect 10892 6244 11144 6272
rect 11284 6244 11620 6272
rect 11844 6272 11900 6300
rect 12936 6272 13104 6300
rect 13160 6328 13356 6356
rect 13664 6328 15092 6356
rect 13160 6272 13384 6328
rect 13636 6300 13916 6328
rect 14028 6300 15120 6328
rect 11844 6244 11928 6272
rect 10332 6216 10752 6244
rect 10920 6216 11172 6244
rect 11312 6216 11648 6244
rect 11872 6216 11928 6244
rect 12936 6216 13132 6272
rect 10332 6188 10724 6216
rect 9772 6160 10276 6188
rect 10304 6160 10724 6188
rect 10920 6188 11200 6216
rect 11312 6188 11676 6216
rect 11872 6188 11956 6216
rect 10920 6160 11228 6188
rect 11340 6160 11704 6188
rect 9520 6132 9576 6160
rect 9604 6132 10696 6160
rect 4592 6104 4760 6132
rect 4564 6076 4760 6104
rect 8036 6104 8484 6132
rect 8596 6104 8848 6132
rect 9184 6104 9268 6132
rect 8036 6076 8456 6104
rect 4564 6048 4732 6076
rect 4536 6020 4732 6048
rect 8008 6048 8456 6076
rect 8568 6076 8820 6104
rect 9240 6076 9324 6104
rect 9408 6076 9464 6132
rect 9548 6104 10696 6132
rect 10892 6104 10948 6160
rect 11004 6132 11256 6160
rect 11368 6132 11704 6160
rect 11900 6132 11956 6188
rect 12964 6160 13132 6216
rect 13188 6244 13384 6272
rect 13608 6272 13832 6300
rect 14084 6272 15148 6300
rect 13608 6244 13804 6272
rect 13916 6244 14000 6272
rect 14112 6244 15148 6272
rect 13188 6160 13412 6244
rect 11032 6104 11284 6132
rect 9548 6076 10668 6104
rect 10864 6076 10920 6104
rect 10948 6076 11284 6104
rect 11396 6076 11732 6132
rect 11900 6104 11984 6132
rect 12964 6104 13160 6160
rect 8568 6048 8792 6076
rect 9268 6048 9352 6076
rect 9436 6048 9464 6076
rect 9492 6048 9828 6076
rect 10192 6048 10668 6076
rect 10836 6048 11004 6076
rect 11088 6048 11312 6076
rect 11424 6048 11760 6076
rect 11928 6048 11984 6104
rect 8008 6020 8428 6048
rect 8540 6020 8764 6048
rect 9324 6020 9408 6048
rect 9436 6020 9716 6048
rect 10248 6020 10640 6048
rect 10780 6020 10920 6048
rect 11088 6020 11340 6048
rect 11424 6020 11788 6048
rect 11928 6020 12012 6048
rect 12992 6020 13160 6104
rect 13216 6132 13412 6160
rect 13580 6216 13636 6244
rect 13664 6216 13776 6244
rect 13860 6216 14056 6244
rect 14140 6216 15064 6244
rect 15092 6216 15176 6244
rect 13580 6160 13608 6216
rect 13692 6188 13776 6216
rect 13832 6188 14084 6216
rect 13692 6160 13748 6188
rect 13580 6132 13748 6160
rect 13216 6048 13440 6132
rect 13608 6048 13748 6132
rect 13244 6020 13440 6048
rect 4536 5992 4704 6020
rect 3668 5880 3836 5908
rect 1904 5824 2072 5852
rect 2520 5824 2688 5852
rect 2996 5824 3164 5852
rect 1876 5712 2072 5824
rect 2492 5712 2688 5824
rect 2968 5712 3164 5824
rect 1876 5684 2044 5712
rect 2492 5684 2660 5712
rect 2968 5684 3136 5712
rect 1848 5572 2044 5684
rect 2464 5600 2660 5684
rect 2940 5600 3136 5684
rect 2464 5572 2632 5600
rect 2940 5572 3108 5600
rect 1848 5544 2016 5572
rect 1820 5432 2016 5544
rect 2436 5460 2632 5572
rect 2912 5460 3108 5572
rect 3276 5516 3444 5852
rect 3640 5768 3836 5880
rect 3612 5656 3808 5768
rect 4200 5712 4368 5992
rect 4508 5964 4704 5992
rect 7980 5992 8428 6020
rect 8512 5992 8764 6020
rect 9352 5992 9632 6020
rect 10220 5992 10640 6020
rect 10696 5992 10864 6020
rect 11116 5992 11340 6020
rect 11452 5992 11788 6020
rect 7980 5964 8400 5992
rect 8512 5964 8792 5992
rect 9352 5964 9576 5992
rect 10220 5964 10752 5992
rect 10808 5964 10836 5992
rect 11144 5964 11368 5992
rect 4508 5936 4676 5964
rect 4480 5908 4676 5936
rect 7952 5908 8372 5964
rect 8484 5936 8708 5964
rect 8764 5936 8820 5964
rect 9324 5936 9520 5964
rect 8484 5908 8680 5936
rect 8792 5908 8848 5936
rect 9296 5908 9492 5936
rect 10192 5908 10696 5964
rect 10780 5936 10836 5964
rect 11172 5936 11368 5964
rect 11480 5936 11816 5992
rect 11956 5936 12012 6020
rect 10780 5908 10808 5936
rect 4480 5880 4648 5908
rect 7952 5880 8344 5908
rect 4452 5852 4648 5880
rect 7924 5852 8344 5880
rect 8456 5880 8680 5908
rect 8456 5852 8652 5880
rect 8820 5852 8876 5908
rect 9268 5880 9436 5908
rect 10164 5880 10724 5908
rect 10752 5880 10808 5908
rect 11172 5880 11396 5936
rect 11508 5880 11844 5936
rect 11956 5908 12040 5936
rect 13020 5908 13188 6020
rect 13244 5936 13468 6020
rect 13636 5992 13748 6048
rect 13804 6020 14112 6188
rect 14168 6160 15036 6216
rect 15120 6160 15176 6216
rect 14168 6132 15176 6160
rect 14168 6020 15148 6132
rect 13832 5992 14084 6020
rect 14168 5992 14336 6020
rect 14728 5992 15148 6020
rect 13664 5964 13776 5992
rect 13860 5964 14084 5992
rect 14140 5964 14336 5992
rect 14392 5964 14700 5992
rect 13664 5936 13804 5964
rect 13888 5936 14028 5964
rect 14140 5936 14364 5964
rect 14392 5936 14672 5964
rect 14728 5936 15120 5992
rect 13272 5908 13468 5936
rect 13692 5908 13832 5936
rect 14084 5908 14364 5936
rect 9240 5852 9408 5880
rect 10164 5852 10556 5880
rect 10584 5852 10780 5880
rect 11032 5852 11424 5880
rect 4452 5796 4620 5852
rect 7924 5824 8316 5852
rect 4424 5740 4592 5796
rect 7896 5768 8316 5824
rect 8428 5824 8652 5852
rect 8848 5824 8904 5852
rect 9212 5824 9380 5852
rect 9912 5824 10080 5852
rect 10136 5824 10780 5852
rect 10864 5824 11116 5852
rect 11228 5824 11424 5852
rect 11536 5824 11872 5880
rect 11984 5824 12040 5908
rect 13048 5824 13216 5908
rect 13272 5824 13496 5908
rect 13692 5880 13860 5908
rect 14056 5880 14392 5908
rect 14420 5880 14644 5936
rect 14700 5908 15120 5936
rect 14700 5880 15092 5908
rect 13720 5852 14392 5880
rect 14448 5852 14616 5880
rect 14672 5852 14952 5880
rect 15008 5852 15092 5880
rect 8428 5796 8624 5824
rect 8876 5796 8932 5824
rect 9184 5796 9352 5824
rect 9772 5796 11060 5824
rect 8400 5768 8624 5796
rect 8904 5768 8960 5796
rect 9156 5768 9324 5796
rect 9716 5768 11060 5796
rect 11256 5768 11452 5824
rect 11564 5796 11900 5824
rect 11984 5796 12068 5824
rect 11564 5768 11928 5796
rect 4200 5684 4340 5712
rect 4424 5684 4564 5740
rect 7896 5712 8288 5768
rect 8400 5740 8652 5768
rect 8932 5740 8988 5768
rect 9156 5740 9296 5768
rect 9660 5740 9940 5768
rect 10052 5740 11088 5768
rect 8372 5712 8680 5740
rect 8932 5712 9016 5740
rect 4200 5656 4536 5684
rect 3612 5628 3780 5656
rect 4200 5628 4508 5656
rect 2436 5432 2604 5460
rect 2912 5432 3080 5460
rect 1792 5320 1988 5432
rect 2408 5320 2604 5432
rect 2884 5320 3080 5432
rect 1792 5292 1960 5320
rect 2408 5292 2576 5320
rect 2884 5292 3052 5320
rect 1764 5180 1960 5292
rect 2380 5208 2576 5292
rect 2856 5208 3052 5292
rect 2380 5180 2548 5208
rect 2856 5180 3024 5208
rect 1764 5152 1932 5180
rect 1736 5040 1932 5152
rect 2352 5068 2548 5180
rect 2828 5068 3024 5180
rect 2352 5040 2520 5068
rect 2828 5040 2996 5068
rect 1736 5012 1904 5040
rect 1708 4928 1904 5012
rect 2324 4928 2520 5040
rect 2800 4928 2996 5040
rect 3304 5040 3444 5516
rect 3584 5516 3780 5628
rect 4228 5600 4508 5628
rect 7868 5628 8260 5712
rect 8372 5656 8568 5712
rect 8652 5684 8708 5712
rect 8960 5684 9016 5712
rect 9128 5684 9268 5740
rect 9604 5712 9828 5740
rect 10080 5712 10472 5740
rect 10528 5712 11088 5740
rect 9576 5684 9744 5712
rect 10080 5684 10444 5712
rect 10584 5684 11088 5712
rect 11284 5712 11480 5768
rect 11564 5740 11956 5768
rect 11592 5712 11984 5740
rect 12012 5712 12068 5796
rect 13076 5712 13244 5824
rect 13300 5796 13496 5824
rect 13748 5824 14420 5852
rect 13748 5796 13832 5824
rect 13888 5796 14420 5824
rect 14476 5824 14616 5852
rect 14644 5824 14924 5852
rect 14476 5796 14588 5824
rect 14644 5796 14952 5824
rect 15008 5796 15064 5852
rect 13300 5712 13524 5796
rect 13776 5768 13804 5796
rect 13888 5768 14448 5796
rect 14504 5768 14588 5796
rect 14616 5768 15064 5796
rect 13776 5740 13832 5768
rect 13888 5740 14476 5768
rect 14504 5740 14560 5768
rect 14616 5740 15036 5768
rect 13804 5712 14476 5740
rect 14588 5712 15036 5740
rect 11284 5684 11508 5712
rect 8680 5656 8736 5684
rect 8988 5656 9044 5684
rect 9100 5656 9240 5684
rect 9548 5656 9688 5684
rect 10052 5656 10444 5684
rect 7868 5600 8232 5628
rect 4228 5544 4480 5600
rect 3584 5488 3752 5516
rect 3556 5376 3752 5488
rect 4228 5488 4452 5544
rect 7840 5516 8232 5600
rect 8344 5600 8540 5656
rect 8708 5628 8764 5656
rect 9016 5628 9212 5656
rect 9520 5628 9660 5656
rect 10052 5628 10472 5656
rect 10612 5628 11060 5684
rect 11312 5656 11508 5684
rect 11592 5656 12068 5712
rect 11284 5628 11508 5656
rect 11620 5628 12068 5656
rect 13104 5684 13244 5712
rect 13328 5684 13524 5712
rect 13832 5684 14504 5712
rect 14560 5684 15008 5712
rect 13104 5628 13272 5684
rect 8736 5600 8820 5628
rect 9044 5600 9212 5628
rect 9492 5600 9632 5628
rect 10024 5600 10500 5628
rect 10584 5600 11032 5628
rect 11228 5600 11536 5628
rect 8344 5572 9184 5600
rect 9464 5572 9576 5600
rect 9856 5572 10528 5600
rect 10556 5572 11060 5600
rect 11200 5572 11284 5600
rect 8316 5544 8540 5572
rect 8792 5544 8904 5572
rect 8988 5544 9184 5572
rect 4228 5404 4424 5488
rect 7840 5460 8204 5516
rect 4228 5376 4396 5404
rect 3528 5264 3724 5376
rect 4200 5264 4396 5376
rect 7812 5348 8204 5460
rect 8316 5488 8512 5544
rect 8848 5516 8904 5544
rect 9044 5516 9156 5544
rect 9436 5516 9548 5572
rect 9800 5544 9884 5572
rect 9996 5544 10388 5572
rect 10444 5544 11060 5572
rect 11144 5544 11228 5572
rect 9744 5516 9800 5544
rect 8876 5488 8932 5516
rect 9016 5488 9156 5516
rect 9408 5488 9520 5516
rect 9716 5488 9772 5516
rect 8316 5432 8484 5488
rect 8904 5460 8960 5488
rect 9016 5460 9128 5488
rect 8932 5432 9128 5460
rect 8288 5348 8484 5432
rect 8960 5404 9128 5432
rect 9380 5432 9492 5488
rect 9688 5460 9772 5488
rect 9996 5488 10360 5544
rect 10472 5516 11172 5544
rect 11340 5516 11536 5600
rect 11620 5600 12096 5628
rect 11620 5572 12012 5600
rect 11648 5544 12012 5572
rect 13132 5572 13272 5628
rect 13328 5600 13552 5684
rect 13832 5656 15008 5684
rect 13860 5628 14980 5656
rect 13860 5600 14952 5628
rect 13356 5572 13552 5600
rect 13888 5572 14952 5600
rect 13132 5544 13300 5572
rect 10472 5488 11144 5516
rect 11340 5488 11564 5516
rect 9996 5460 10388 5488
rect 10472 5460 11172 5488
rect 9660 5432 9800 5460
rect 10024 5432 11200 5460
rect 9380 5404 9464 5432
rect 9632 5404 9688 5432
rect 9744 5404 9828 5432
rect 8876 5376 9100 5404
rect 8596 5348 9100 5376
rect 3528 5236 3696 5264
rect 4200 5236 4368 5264
rect 3500 5124 3696 5236
rect 4172 5124 4368 5236
rect 3500 5068 3668 5124
rect 4172 5096 4340 5124
rect 3472 5040 3668 5068
rect 3304 4984 3668 5040
rect 4144 4984 4340 5096
rect 1708 4900 1876 4928
rect 2324 4900 2492 4928
rect 2800 4900 2968 4928
rect 1680 4788 1876 4900
rect 2296 4788 2492 4900
rect 2772 4788 2968 4900
rect 3304 4844 3640 4984
rect 4116 4872 4312 4984
rect 7812 4900 8176 5348
rect 8288 5320 8708 5348
rect 8288 5292 8484 5320
rect 8288 5012 8456 5292
rect 8988 5264 9100 5348
rect 9352 5376 9464 5404
rect 9604 5376 9660 5404
rect 9772 5376 9856 5404
rect 10052 5376 11200 5432
rect 11368 5404 11564 5488
rect 11648 5460 12040 5544
rect 13160 5460 13300 5544
rect 13356 5516 13580 5572
rect 13916 5544 14924 5572
rect 13384 5488 13580 5516
rect 13944 5516 14728 5544
rect 14784 5516 14896 5544
rect 13944 5488 14084 5516
rect 14112 5488 14700 5516
rect 14812 5488 14868 5516
rect 11340 5376 11564 5404
rect 9352 5320 9436 5376
rect 9604 5348 9632 5376
rect 9800 5348 9884 5376
rect 8960 5236 9100 5264
rect 9324 5292 9436 5320
rect 9576 5320 9632 5348
rect 9828 5320 9912 5348
rect 10052 5320 10108 5376
rect 10136 5348 10248 5376
rect 10304 5348 11200 5376
rect 11284 5348 11564 5376
rect 11676 5348 12040 5460
rect 13188 5404 13328 5460
rect 13384 5404 13608 5488
rect 13972 5460 14056 5488
rect 14000 5432 14056 5460
rect 14140 5460 14728 5488
rect 14784 5460 14868 5488
rect 14140 5432 14840 5460
rect 14028 5404 14812 5432
rect 13216 5348 13328 5404
rect 13412 5376 13608 5404
rect 14056 5376 14784 5404
rect 10360 5320 11172 5348
rect 11228 5320 11312 5348
rect 8960 5096 9072 5236
rect 8960 5068 9100 5096
rect 8288 4984 8596 5012
rect 8288 4956 8736 4984
rect 8988 4956 9100 5068
rect 9324 5040 9408 5292
rect 9576 5236 9604 5320
rect 9856 5292 10108 5320
rect 9884 5264 10108 5292
rect 9884 5236 9968 5264
rect 10024 5236 10108 5264
rect 10388 5292 11256 5320
rect 10388 5236 11200 5292
rect 11396 5236 11592 5348
rect 11676 5236 12068 5348
rect 13216 5320 13356 5348
rect 13244 5236 13356 5320
rect 13412 5320 13636 5376
rect 13664 5348 13804 5376
rect 14084 5348 14756 5376
rect 13664 5320 13692 5348
rect 13804 5320 13860 5348
rect 14112 5320 14700 5348
rect 13412 5292 13664 5320
rect 13860 5292 13944 5320
rect 14140 5292 14672 5320
rect 9548 5208 9604 5236
rect 9548 5124 9576 5208
rect 9856 5124 9912 5236
rect 10080 5208 10136 5236
rect 10080 5180 10164 5208
rect 10388 5180 11116 5236
rect 11144 5208 11312 5236
rect 11424 5208 11592 5236
rect 11256 5180 11592 5208
rect 10080 5152 10332 5180
rect 10388 5152 11144 5180
rect 11368 5152 11592 5180
rect 10080 5124 11172 5152
rect 9548 5096 9604 5124
rect 9856 5096 9940 5124
rect 10080 5096 10136 5124
rect 10360 5096 11172 5124
rect 9324 5012 9436 5040
rect 9352 4956 9436 5012
rect 9576 5012 9604 5096
rect 9828 5068 9968 5096
rect 10024 5068 10108 5096
rect 9772 5040 10108 5068
rect 10388 5068 10444 5096
rect 10472 5068 11172 5096
rect 9744 5012 9856 5040
rect 9968 5012 10080 5040
rect 10388 5012 10416 5068
rect 10500 5040 11172 5068
rect 9576 4984 9632 5012
rect 9688 4984 9800 5012
rect 9604 4956 9744 4984
rect 4116 4844 4284 4872
rect 1680 4760 1848 4788
rect 1652 4704 1848 4760
rect 2268 4704 2464 4788
rect 2744 4704 2940 4788
rect 3304 4732 3612 4844
rect 4088 4732 4284 4844
rect 7812 4788 8204 4900
rect 8288 4844 8484 4956
rect 8596 4928 8876 4956
rect 8988 4928 9128 4956
rect 9352 4928 9464 4956
rect 9604 4928 9688 4956
rect 8736 4900 9128 4928
rect 8876 4872 9128 4900
rect 9380 4900 9464 4928
rect 9632 4900 9688 4928
rect 9380 4872 9492 4900
rect 9660 4872 9716 4900
rect 10052 4872 10108 5012
rect 10360 4984 10416 5012
rect 10556 5012 11172 5040
rect 11424 5012 11592 5152
rect 11704 5012 12068 5236
rect 13272 5180 13384 5236
rect 13440 5180 13664 5292
rect 13916 5264 14000 5292
rect 14168 5264 14336 5292
rect 14000 5236 14056 5264
rect 14196 5236 14336 5264
rect 14420 5264 14644 5292
rect 14420 5236 14588 5264
rect 14056 5208 14112 5236
rect 14252 5208 14532 5236
rect 14112 5180 14168 5208
rect 14280 5180 14476 5208
rect 13300 5124 13384 5180
rect 13468 5152 13664 5180
rect 14168 5152 14252 5180
rect 14336 5152 14420 5180
rect 13300 5096 13412 5124
rect 13328 5040 13412 5096
rect 13468 5068 13692 5152
rect 14252 5124 14336 5152
rect 13916 5096 13944 5124
rect 14084 5096 14112 5124
rect 14224 5096 14252 5124
rect 14336 5096 14476 5124
rect 13496 5040 13720 5068
rect 13888 5040 13972 5096
rect 14056 5068 14140 5096
rect 14056 5040 14112 5068
rect 14196 5040 14280 5096
rect 14448 5068 14728 5096
rect 14728 5040 14784 5068
rect 13328 5012 13440 5040
rect 13496 5012 13748 5040
rect 14784 5012 14812 5040
rect 10556 4984 11200 5012
rect 10360 4956 10388 4984
rect 10556 4956 10640 4984
rect 10696 4956 11088 4984
rect 11144 4956 11256 4984
rect 10332 4928 10388 4956
rect 10304 4900 10360 4928
rect 10528 4900 10640 4956
rect 10892 4928 11004 4956
rect 11228 4928 11312 4956
rect 10276 4872 10332 4900
rect 8988 4844 9128 4872
rect 9408 4844 9492 4872
rect 9688 4844 9744 4872
rect 8288 4816 8512 4844
rect 8988 4816 9156 4844
rect 9408 4816 9520 4844
rect 9716 4816 9772 4844
rect 7840 4760 8204 4788
rect 3304 4704 3584 4732
rect 4088 4704 4256 4732
rect 7840 4648 8232 4760
rect 8316 4732 8512 4816
rect 8960 4788 9156 4816
rect 9436 4788 9548 4816
rect 9744 4788 9828 4816
rect 10080 4788 10136 4872
rect 10248 4844 10304 4872
rect 10500 4844 10612 4900
rect 10864 4872 11004 4928
rect 11284 4900 11368 4928
rect 11396 4900 11592 5012
rect 11676 4900 12068 5012
rect 13356 4956 13440 5012
rect 13524 4984 13776 5012
rect 13524 4956 13804 4984
rect 13972 4956 14056 5012
rect 14140 4956 14224 5012
rect 14308 4984 14364 5012
rect 14812 4984 14840 5012
rect 14280 4956 14364 4984
rect 14840 4956 14868 4984
rect 13356 4928 13468 4956
rect 13384 4900 13468 4928
rect 13552 4928 13860 4956
rect 14000 4928 14028 4956
rect 14168 4928 14196 4956
rect 14308 4928 14336 4956
rect 14840 4928 14896 4956
rect 13552 4900 13944 4928
rect 14840 4900 14924 4928
rect 11340 4872 11564 4900
rect 10864 4844 10976 4872
rect 10220 4816 10276 4844
rect 10472 4816 10584 4844
rect 10164 4788 10248 4816
rect 8932 4760 9016 4788
rect 9044 4760 9184 4788
rect 9436 4760 9576 4788
rect 9800 4760 9884 4788
rect 10080 4760 10192 4788
rect 10444 4760 10556 4816
rect 10836 4788 10976 4844
rect 11396 4816 11564 4872
rect 11676 4816 12040 4900
rect 13412 4872 13468 4900
rect 13580 4872 15484 4900
rect 13412 4844 13496 4872
rect 13608 4844 15484 4872
rect 13440 4816 13524 4844
rect 13636 4816 15484 4844
rect 8876 4732 9184 4760
rect 9464 4732 9604 4760
rect 9856 4732 10136 4760
rect 10416 4732 10528 4760
rect 10808 4732 10948 4788
rect 11368 4732 11564 4816
rect 8316 4704 8540 4732
rect 8568 4704 9212 4732
rect 9492 4704 9632 4732
rect 10388 4704 10500 4732
rect 10780 4704 10920 4732
rect 11368 4704 11536 4732
rect 8344 4676 8932 4704
rect 9072 4676 9212 4704
rect 9520 4676 9660 4704
rect 10332 4676 10472 4704
rect 10780 4676 11116 4704
rect 11340 4676 11536 4704
rect 11648 4704 12040 4816
rect 13468 4788 13552 4816
rect 13664 4788 15484 4816
rect 13468 4760 13580 4788
rect 13720 4760 15484 4788
rect 13496 4732 13608 4760
rect 13776 4732 15484 4760
rect 13524 4704 13636 4732
rect 13860 4704 15484 4732
rect 11648 4676 12012 4704
rect 13552 4676 13692 4704
rect 7868 4564 8260 4648
rect 8344 4592 8540 4676
rect 8820 4648 8904 4676
rect 9100 4648 9240 4676
rect 9548 4648 9688 4676
rect 10304 4648 10444 4676
rect 10752 4648 10920 4676
rect 11032 4648 11536 4676
rect 8792 4620 8876 4648
rect 9100 4620 9268 4648
rect 9576 4620 9744 4648
rect 10248 4620 10416 4648
rect 10724 4620 10920 4648
rect 8764 4592 8848 4620
rect 9072 4592 9268 4620
rect 9604 4592 9828 4620
rect 10164 4592 10388 4620
rect 10724 4592 10864 4620
rect 10892 4592 10948 4620
rect 7868 4536 8288 4564
rect 7896 4480 8288 4536
rect 8372 4536 8568 4592
rect 8736 4564 8820 4592
rect 9044 4564 9128 4592
rect 9156 4564 9296 4592
rect 9660 4564 9968 4592
rect 10024 4564 10332 4592
rect 10696 4564 10836 4592
rect 10920 4564 10976 4592
rect 11312 4564 11508 4648
rect 11620 4592 12012 4676
rect 13608 4648 13776 4676
rect 13636 4620 13888 4648
rect 13692 4592 15260 4620
rect 8708 4536 8792 4564
rect 9016 4536 9100 4564
rect 9184 4536 9324 4564
rect 9716 4536 10276 4564
rect 10668 4536 10836 4564
rect 8372 4508 8596 4536
rect 8680 4508 8764 4536
rect 8988 4508 9072 4536
rect 9184 4508 9352 4536
rect 9800 4508 10220 4536
rect 10640 4508 10864 4536
rect 10948 4508 11004 4564
rect 11284 4508 11480 4564
rect 11592 4508 11984 4592
rect 13776 4564 15260 4592
rect 8400 4480 8596 4508
rect 8652 4480 8736 4508
rect 8960 4480 9044 4508
rect 9212 4480 9380 4508
rect 9940 4480 10052 4508
rect 10612 4480 11032 4508
rect 11256 4480 11480 4508
rect 11564 4480 11984 4508
rect 7896 4452 8316 4480
rect 8400 4452 8708 4480
rect 8932 4452 9016 4480
rect 9240 4452 9408 4480
rect 10584 4452 10808 4480
rect 10920 4452 11144 4480
rect 11256 4452 11452 4480
rect 11564 4452 11956 4480
rect 7924 4424 8316 4452
rect 8428 4424 8680 4452
rect 8932 4424 8988 4452
rect 9268 4424 9464 4452
rect 10556 4424 10724 4452
rect 2744 4396 3500 4424
rect 4648 4396 4900 4424
rect 5572 4396 5824 4424
rect 6412 4396 6664 4424
rect 7028 4396 7252 4424
rect 2856 4368 3780 4396
rect 4004 4368 4172 4396
rect 4704 4368 5236 4396
rect 5600 4368 6216 4396
rect 6440 4368 6804 4396
rect 7084 4368 7392 4396
rect 7924 4368 8344 4424
rect 8428 4396 8652 4424
rect 8904 4396 8960 4424
rect 9296 4396 9492 4424
rect 10500 4396 10696 4424
rect 10780 4396 10836 4452
rect 11032 4424 11452 4452
rect 11060 4396 11116 4424
rect 3192 4284 3780 4368
rect 3192 4228 3752 4284
rect 3976 4256 4172 4368
rect 4872 4340 5236 4368
rect 5768 4340 6244 4368
rect 4900 4312 5236 4340
rect 5740 4312 6244 4340
rect 3976 4228 4144 4256
rect 4872 4228 5236 4312
rect 5712 4284 6272 4312
rect 5684 4256 6300 4284
rect 6608 4256 6804 4368
rect 7196 4340 7392 4368
rect 7952 4340 8344 4368
rect 8456 4368 8652 4396
rect 8876 4368 8960 4396
rect 9324 4368 9548 4396
rect 10472 4368 10668 4396
rect 10808 4368 10864 4396
rect 11060 4368 11144 4396
rect 8456 4340 8680 4368
rect 8848 4340 8932 4368
rect 9352 4340 9576 4368
rect 10416 4340 10640 4368
rect 10836 4340 10864 4368
rect 11088 4340 11144 4368
rect 11200 4368 11424 4424
rect 11536 4396 11956 4452
rect 11536 4368 11928 4396
rect 11200 4340 11396 4368
rect 7196 4312 7364 4340
rect 5628 4228 6328 4256
rect 6608 4228 6776 4256
rect 3164 4116 3360 4228
rect 3948 4116 4144 4228
rect 4844 4172 5012 4228
rect 5040 4200 5236 4228
rect 4844 4144 4984 4172
rect 5068 4144 5236 4200
rect 5600 4200 5880 4228
rect 6076 4200 6356 4228
rect 5600 4172 5852 4200
rect 6104 4172 6356 4200
rect 5600 4144 5824 4172
rect 6104 4144 6328 4172
rect 3164 4088 3332 4116
rect 3948 4088 4116 4116
rect 4816 4088 4984 4144
rect 3136 3976 3332 4088
rect 3920 3976 4116 4088
rect 4788 4060 4984 4088
rect 4788 4004 4956 4060
rect 4760 3976 4956 4004
rect 3108 3864 3304 3976
rect 3892 3864 4088 3976
rect 4760 3920 4928 3976
rect 4732 3892 4928 3920
rect 5040 3892 5208 4144
rect 5572 4060 5768 4144
rect 5572 4032 5740 4060
rect 5544 3920 5740 4032
rect 6132 4032 6328 4144
rect 6580 4116 6776 4228
rect 7168 4200 7364 4312
rect 7952 4312 8372 4340
rect 8484 4312 8680 4340
rect 8820 4312 8904 4340
rect 9408 4312 9660 4340
rect 10332 4312 10584 4340
rect 10836 4312 10892 4340
rect 11116 4312 11396 4340
rect 11508 4312 11928 4368
rect 7952 4284 8400 4312
rect 8484 4284 8708 4312
rect 8792 4284 8876 4312
rect 9436 4284 9716 4312
rect 10276 4284 10556 4312
rect 10864 4284 10892 4312
rect 7980 4256 8400 4284
rect 8512 4256 8736 4284
rect 8764 4256 8848 4284
rect 9408 4256 9828 4284
rect 10164 4256 10500 4284
rect 10864 4256 10920 4284
rect 11144 4256 11368 4312
rect 11480 4284 11900 4312
rect 11452 4256 11900 4284
rect 7980 4228 8428 4256
rect 8512 4228 8820 4256
rect 9352 4228 9464 4256
rect 9492 4228 10444 4256
rect 8008 4200 8428 4228
rect 8540 4200 8792 4228
rect 9296 4200 9408 4228
rect 7168 4172 7336 4200
rect 8008 4172 8456 4200
rect 8568 4172 8792 4200
rect 9240 4172 9352 4200
rect 9492 4172 9548 4228
rect 9604 4200 10444 4228
rect 10892 4200 10948 4256
rect 11116 4228 11340 4256
rect 11452 4228 11872 4256
rect 11088 4200 11312 4228
rect 9576 4172 10304 4200
rect 10332 4172 10472 4200
rect 10920 4172 10976 4200
rect 6580 4088 6748 4116
rect 6132 4004 6300 4032
rect 5544 3892 5712 3920
rect 3108 3836 3276 3864
rect 3892 3836 4060 3864
rect 4732 3836 4900 3892
rect 3080 3724 3276 3836
rect 3864 3724 4060 3836
rect 4704 3808 4900 3836
rect 4704 3780 4872 3808
rect 4676 3724 4872 3780
rect 3080 3696 3248 3724
rect 3864 3696 4032 3724
rect 4676 3696 4844 3724
rect 3052 3584 3248 3696
rect 3836 3584 4032 3696
rect 4648 3668 4844 3696
rect 5012 3668 5208 3892
rect 5516 3780 5712 3892
rect 6104 3892 6300 4004
rect 6552 3976 6748 4088
rect 7140 4060 7336 4172
rect 8036 4116 8484 4172
rect 8568 4144 8820 4172
rect 9212 4144 9324 4172
rect 9492 4144 9632 4172
rect 8596 4116 8848 4144
rect 9156 4116 9268 4144
rect 9492 4116 9604 4144
rect 8064 4088 8512 4116
rect 8624 4088 8876 4116
rect 9100 4088 9212 4116
rect 9492 4088 9576 4116
rect 8064 4060 8540 4088
rect 8652 4060 8904 4088
rect 9044 4060 9156 4088
rect 9464 4060 9548 4088
rect 7140 4032 7308 4060
rect 8092 4032 8540 4060
rect 8680 4032 8932 4060
rect 8988 4032 9100 4060
rect 9408 4032 9548 4060
rect 9660 4032 9716 4172
rect 9800 4144 10248 4172
rect 10136 4116 10276 4144
rect 6104 3864 6272 3892
rect 6076 3836 6272 3864
rect 6524 3864 6720 3976
rect 7112 3948 7308 4032
rect 8120 4004 8568 4032
rect 8680 4004 9072 4032
rect 9380 4004 9548 4032
rect 8120 3976 8596 4004
rect 8708 3976 9016 4004
rect 9352 3976 9436 4004
rect 8148 3948 8624 3976
rect 8736 3948 9016 3976
rect 9324 3948 9408 3976
rect 9492 3948 9520 4004
rect 7112 3892 7280 3948
rect 8148 3920 8652 3948
rect 8764 3920 9072 3948
rect 9296 3920 9380 3948
rect 8176 3892 8680 3920
rect 8792 3892 9100 3920
rect 9268 3892 9352 3920
rect 6524 3836 6692 3864
rect 5516 3752 5740 3780
rect 5488 3724 5768 3752
rect 6496 3724 6692 3836
rect 7084 3808 7280 3892
rect 8204 3864 8708 3892
rect 8848 3864 9156 3892
rect 9240 3864 9324 3892
rect 8232 3836 8736 3864
rect 8876 3836 9296 3864
rect 8232 3808 8764 3836
rect 8904 3808 9268 3836
rect 7084 3780 7252 3808
rect 8260 3780 8792 3808
rect 8932 3780 9296 3808
rect 5488 3696 5796 3724
rect 6496 3696 6664 3724
rect 5516 3668 5824 3696
rect 4648 3612 4816 3668
rect 4620 3584 4816 3612
rect 3052 3556 3584 3584
rect 3836 3556 4004 3584
rect 3024 3528 3584 3556
rect 3024 3444 3556 3528
rect 3808 3472 4004 3556
rect 4620 3528 4788 3584
rect 4592 3500 4788 3528
rect 5012 3500 5180 3668
rect 5544 3640 5852 3668
rect 5572 3612 5880 3640
rect 5600 3584 5908 3612
rect 6468 3584 6664 3696
rect 7056 3668 7252 3780
rect 8288 3752 8820 3780
rect 8988 3752 9352 3780
rect 8316 3724 8848 3752
rect 9016 3724 9436 3752
rect 9464 3724 9520 3948
rect 8344 3696 8904 3724
rect 9072 3696 9520 3724
rect 9688 3920 9716 4032
rect 10108 4088 10192 4116
rect 10220 4088 10304 4116
rect 10108 4004 10164 4088
rect 10248 4060 10304 4088
rect 10332 4060 10388 4172
rect 10416 4144 10500 4172
rect 10948 4144 10976 4172
rect 11060 4172 11312 4200
rect 11424 4200 11872 4228
rect 11424 4172 11844 4200
rect 11060 4144 11284 4172
rect 11396 4144 11844 4172
rect 10444 4116 10528 4144
rect 10948 4116 11004 4144
rect 11032 4116 11256 4144
rect 10472 4088 10556 4116
rect 10976 4088 11256 4116
rect 11368 4088 11816 4144
rect 10500 4060 10584 4088
rect 10976 4060 11228 4088
rect 11340 4060 11788 4088
rect 10248 4032 10388 4060
rect 10528 4032 10584 4060
rect 10948 4032 11200 4060
rect 11312 4032 11788 4060
rect 10276 4004 10360 4032
rect 10528 4004 10612 4032
rect 10920 4004 11172 4032
rect 11284 4004 11760 4032
rect 10080 3920 10136 4004
rect 8372 3668 8932 3696
rect 9100 3668 9604 3696
rect 9688 3668 9744 3920
rect 10052 3892 10136 3920
rect 10304 3976 10360 4004
rect 10556 3976 10640 4004
rect 10864 3976 11144 4004
rect 11284 3976 11732 4004
rect 10304 3920 10388 3976
rect 10584 3948 10668 3976
rect 10836 3948 11116 3976
rect 11256 3948 11732 3976
rect 10612 3920 10696 3948
rect 10808 3920 11088 3948
rect 11228 3920 11704 3948
rect 10304 3892 10416 3920
rect 10640 3892 10696 3920
rect 10752 3892 11060 3920
rect 11200 3892 11676 3920
rect 10052 3808 10108 3892
rect 10304 3864 10444 3892
rect 10304 3808 10360 3864
rect 10388 3836 10444 3864
rect 10668 3864 11032 3892
rect 11172 3864 11676 3892
rect 10668 3836 11004 3864
rect 11144 3836 11648 3864
rect 10416 3808 10472 3836
rect 10640 3808 10976 3836
rect 11116 3808 11620 3836
rect 10024 3724 10080 3808
rect 10304 3780 10332 3808
rect 10416 3780 10500 3808
rect 10584 3780 10920 3808
rect 11088 3780 11592 3808
rect 7056 3640 7224 3668
rect 8372 3640 8988 3668
rect 9156 3640 9772 3668
rect 9996 3640 10052 3724
rect 10276 3696 10332 3780
rect 10444 3752 10892 3780
rect 11032 3752 11592 3780
rect 10444 3724 10836 3752
rect 11004 3724 11564 3752
rect 10360 3696 10808 3724
rect 10976 3696 11536 3724
rect 10248 3668 10752 3696
rect 10920 3668 11508 3696
rect 10080 3640 10696 3668
rect 10892 3640 11480 3668
rect 7028 3584 7224 3640
rect 8400 3612 9016 3640
rect 9212 3612 10640 3640
rect 10836 3612 11452 3640
rect 8428 3584 9072 3612
rect 9268 3584 10584 3612
rect 10808 3584 11424 3612
rect 5628 3556 5936 3584
rect 6468 3556 7224 3584
rect 8484 3556 9128 3584
rect 9352 3556 10528 3584
rect 10752 3556 11396 3584
rect 5656 3528 5936 3556
rect 6440 3528 7224 3556
rect 8512 3528 9184 3556
rect 9436 3528 10444 3556
rect 10696 3528 11368 3556
rect 4592 3472 4760 3500
rect 3808 3444 3976 3472
rect 2996 3416 3556 3444
rect 2996 3332 3192 3416
rect 3780 3332 3976 3444
rect 4564 3416 4760 3472
rect 4564 3388 4732 3416
rect 4536 3332 4732 3388
rect 2996 3304 3164 3332
rect 3780 3304 3948 3332
rect 4536 3304 4704 3332
rect 2968 3192 3164 3304
rect 3752 3192 3948 3304
rect 4508 3276 4704 3304
rect 4508 3248 4676 3276
rect 4984 3248 5180 3500
rect 5684 3500 5964 3528
rect 5684 3472 5992 3500
rect 5712 3444 6020 3472
rect 6440 3444 7196 3528
rect 8540 3500 9240 3528
rect 9520 3500 10332 3528
rect 10640 3500 11340 3528
rect 8568 3472 9296 3500
rect 9688 3472 10192 3500
rect 10556 3472 11312 3500
rect 8596 3444 9380 3472
rect 10472 3444 11256 3472
rect 5740 3416 6048 3444
rect 6412 3416 7196 3444
rect 8624 3416 9492 3444
rect 10388 3416 11228 3444
rect 5768 3388 6076 3416
rect 5796 3360 6104 3388
rect 5824 3332 6132 3360
rect 6412 3332 6608 3416
rect 7000 3388 7168 3416
rect 8680 3388 9604 3416
rect 10276 3388 11200 3416
rect 5852 3304 6160 3332
rect 6412 3304 6580 3332
rect 5880 3276 6160 3304
rect 5908 3248 6160 3276
rect 4508 3220 5180 3248
rect 4480 3192 5180 3220
rect 5936 3220 6160 3248
rect 2968 3164 3136 3192
rect 3752 3164 3920 3192
rect 4480 3164 5152 3192
rect 5236 3164 5572 3192
rect 2940 3052 3136 3164
rect 3724 3052 3920 3164
rect 4452 3080 5152 3164
rect 5376 3108 5572 3164
rect 2912 2940 3108 3052
rect 3696 2940 3892 3052
rect 4424 3024 4620 3080
rect 4424 2996 4592 3024
rect 4396 2940 4592 2996
rect 2912 2912 3080 2940
rect 3696 2912 3864 2940
rect 2884 2800 3080 2912
rect 3668 2800 3864 2912
rect 4368 2856 4564 2940
rect 2884 2772 3052 2800
rect 3668 2772 3836 2800
rect 4340 2772 4536 2856
rect 2856 2660 3052 2772
rect 3640 2744 3836 2772
rect 3640 2688 4200 2744
rect 4312 2716 4508 2772
rect 4956 2744 5152 3080
rect 5348 2996 5544 3108
rect 5936 3080 6132 3220
rect 6384 3192 6580 3304
rect 6972 3276 7168 3388
rect 8708 3360 9800 3388
rect 10080 3360 11144 3388
rect 8764 3332 11116 3360
rect 8792 3304 11060 3332
rect 8848 3276 11032 3304
rect 6972 3248 7140 3276
rect 8904 3248 10976 3276
rect 6384 3164 6552 3192
rect 5348 2968 5516 2996
rect 5320 2884 5516 2968
rect 5908 2968 6104 3080
rect 6356 3052 6552 3164
rect 6944 3136 7140 3248
rect 8932 3220 10920 3248
rect 8988 3192 10864 3220
rect 9072 3164 10808 3192
rect 9128 3136 10752 3164
rect 6944 3108 7112 3136
rect 9184 3108 10668 3136
rect 5908 2940 6076 2968
rect 5320 2856 5488 2884
rect 5880 2856 6076 2940
rect 6328 2940 6524 3052
rect 6916 3024 7112 3108
rect 9268 3080 10584 3108
rect 9380 3052 10500 3080
rect 9492 3024 10360 3052
rect 6916 2996 7084 3024
rect 9660 2996 10192 3024
rect 6328 2912 6496 2940
rect 5292 2800 5516 2856
rect 5852 2828 6076 2856
rect 5824 2800 6048 2828
rect 5292 2772 5544 2800
rect 5796 2772 6048 2800
rect 6300 2800 6496 2912
rect 6888 2884 7084 2996
rect 6888 2856 7056 2884
rect 6300 2772 6468 2800
rect 5292 2744 5572 2772
rect 5768 2744 6048 2772
rect 4928 2716 5152 2744
rect 5320 2716 5992 2744
rect 4312 2688 4480 2716
rect 3640 2660 4172 2688
rect 2828 2576 3024 2660
rect 3612 2576 4172 2660
rect 4284 2632 4480 2688
rect 4256 2576 4452 2632
rect 4928 2576 5124 2716
rect 5348 2688 5964 2716
rect 5376 2660 5936 2688
rect 6272 2660 6468 2772
rect 6860 2744 7056 2856
rect 6860 2716 7028 2744
rect 5376 2632 5908 2660
rect 5404 2604 5852 2632
rect 5432 2576 5824 2604
rect 6244 2576 6440 2660
rect 6832 2632 7028 2716
rect 6832 2604 7000 2632
rect 6804 2576 7000 2604
<< end >>
