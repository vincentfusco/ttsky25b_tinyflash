* SPICE3 file created from tt_um_tinychaos.ext - technology: sky130A

X0 flashADC_3bit_0/vbias_generation_0/XR_bias_2/R2 flashADC_3bit_0/comp_p_6/vbias_p VGND sky130_fd_pr__res_xhigh_po_1p41 l=7
X1 flashADC_3bit_0/vbias_generation_0/XR_bias_3/R2 flashADC_3bit_0/vbias_generation_0/XR_bias_2/R2 VGND sky130_fd_pr__res_xhigh_po_1p41 l=7
X2 flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 flashADC_3bit_0/vbias_generation_0/XR_bias_3/R2 VGND sky130_fd_pr__res_xhigh_po_1p41 l=7
X3 flashADC_3bit_0/vbias_generation_0/XR_bias_4/R1 flashADC_3bit_0/vbias_generation_0/bias_n VGND sky130_fd_pr__res_xhigh_po_1p41 l=7
X4 VGND flashADC_3bit_0/vbias_generation_0/bias_n flashADC_3bit_0/vbias_generation_0/bias_n VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X5 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_6/vbias_p VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X6 flashADC_3bit_0/comp_p_6/vinn ua[1] VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X7 flashADC_3bit_0/comp_p_6/vinn ua[1] VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X8 flashADC_3bit_0/comp_p_1/vinn VGND VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X9 flashADC_3bit_0/comp_p_6/vinn flashADC_3bit_0/comp_p_5/vinn VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X10 flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_5/vinn VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X11 flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_3/vinn VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X12 flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_3/vinn VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X13 flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_0/vinn VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X14 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_0/vinn VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X15 flashADC_3bit_0/comp_p_1/vinn VGND VGND sky130_fd_pr__res_xhigh_po_5p73 l=5.73
X16 flashADC_3bit_0/comp_p_1/latch_right flashADC_3bit_0/comp_p_1/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
X17 VDPWR flashADC_3bit_0/comp_p_1/out_left uo_out[3] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
X18 flashADC_3bit_0/comp_p_1/latch_left flashADC_3bit_0/comp_p_1/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X19 flashADC_3bit_0/comp_p_1/latch_left flashADC_3bit_0/comp_p_1/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=65.25 ps=488.86 w=5 l=1
X20 flashADC_3bit_0/comp_p_1/latch_right flashADC_3bit_0/comp_p_1/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=4 l=1
X21 VDPWR flashADC_3bit_0/comp_p_1/out_left flashADC_3bit_0/comp_p_1/out_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=69.6 pd=506.68 as=2.32 ps=16.58 w=8 l=1
X22 flashADC_3bit_0/comp_p_1/out_left flashADC_3bit_0/comp_p_1/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X23 uo_out[3] flashADC_3bit_0/comp_p_1/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X24 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_1/tail VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X25 flashADC_3bit_0/comp_p_1/tail flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_1/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X26 flashADC_3bit_0/comp_p_1/tail ua[0] flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X27 flashADC_3bit_0/comp_p_1/tail ua[0] flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X28 flashADC_3bit_0/comp_p_1/tail ua[0] flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X29 flashADC_3bit_0/comp_p_1/tail ua[0] flashADC_3bit_0/comp_p_1/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X30 flashADC_3bit_0/comp_p_1/tail flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_1/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X31 flashADC_3bit_0/comp_p_1/tail flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_1/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X32 flashADC_3bit_0/comp_p_1/tail flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_1/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X33 flashADC_3bit_0/comp_p_0/latch_right flashADC_3bit_0/comp_p_0/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=5 l=1
X34 VDPWR flashADC_3bit_0/comp_p_0/out_left uo_out[4] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X35 flashADC_3bit_0/comp_p_0/latch_left flashADC_3bit_0/comp_p_0/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=4 l=1
X36 flashADC_3bit_0/comp_p_0/latch_left flashADC_3bit_0/comp_p_0/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=5 l=1
X37 flashADC_3bit_0/comp_p_0/latch_right flashADC_3bit_0/comp_p_0/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
X38 VDPWR flashADC_3bit_0/comp_p_0/out_left flashADC_3bit_0/comp_p_0/out_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X39 flashADC_3bit_0/comp_p_0/out_left flashADC_3bit_0/comp_p_0/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X40 uo_out[4] flashADC_3bit_0/comp_p_0/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X41 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_0/tail VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=20.433426 ps=144.985 w=10 l=1
X42 flashADC_3bit_0/comp_p_0/tail flashADC_3bit_0/comp_p_0/vinn flashADC_3bit_0/comp_p_0/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.5942 ps=82.28 w=9.995 l=0.35
X43 flashADC_3bit_0/comp_p_0/tail ua[0] flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.295525 ps=79.645 w=9.995 l=0.35
X44 flashADC_3bit_0/comp_p_0/tail ua[0] flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X45 flashADC_3bit_0/comp_p_0/tail ua[0] flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X46 flashADC_3bit_0/comp_p_0/tail ua[0] flashADC_3bit_0/comp_p_0/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X47 flashADC_3bit_0/comp_p_0/tail flashADC_3bit_0/comp_p_0/vinn flashADC_3bit_0/comp_p_0/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X48 flashADC_3bit_0/comp_p_0/tail flashADC_3bit_0/comp_p_0/vinn flashADC_3bit_0/comp_p_0/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X49 flashADC_3bit_0/comp_p_0/tail flashADC_3bit_0/comp_p_0/vinn flashADC_3bit_0/comp_p_0/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X50 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_2/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=5 l=1
X51 VDPWR flashADC_3bit_0/comp_p_2/out_left uo_out[5] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X52 flashADC_3bit_0/comp_p_2/latch_left flashADC_3bit_0/comp_p_2/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=4 l=1
X53 flashADC_3bit_0/comp_p_2/latch_left flashADC_3bit_0/comp_p_2/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=5 l=1
X54 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_2/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
X55 VDPWR flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/comp_p_2/out_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X56 flashADC_3bit_0/comp_p_2/out_left flashADC_3bit_0/comp_p_2/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X57 uo_out[5] flashADC_3bit_0/comp_p_2/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X58 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_2/tail VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=20.433426 ps=144.985 w=10 l=1
X59 flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_2/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.5942 ps=82.28 w=9.995 l=0.35
X60 flashADC_3bit_0/comp_p_2/tail ua[0] flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.295525 ps=79.645 w=9.995 l=0.35
X61 flashADC_3bit_0/comp_p_2/tail ua[0] flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X62 flashADC_3bit_0/comp_p_2/tail ua[0] flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X63 flashADC_3bit_0/comp_p_2/tail ua[0] flashADC_3bit_0/comp_p_2/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X64 flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_2/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X65 flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_2/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X66 flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_2/vinn flashADC_3bit_0/comp_p_2/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X67 flashADC_3bit_0/comp_p_3/latch_right flashADC_3bit_0/comp_p_3/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=5 l=1
X68 VDPWR flashADC_3bit_0/comp_p_3/out_left uo_out[6] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X69 flashADC_3bit_0/comp_p_3/latch_left flashADC_3bit_0/comp_p_3/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=4 l=1
X70 flashADC_3bit_0/comp_p_3/latch_left flashADC_3bit_0/comp_p_3/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=5 l=1
X71 flashADC_3bit_0/comp_p_3/latch_right flashADC_3bit_0/comp_p_3/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
X72 VDPWR flashADC_3bit_0/comp_p_3/out_left flashADC_3bit_0/comp_p_3/out_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X73 flashADC_3bit_0/comp_p_3/out_left flashADC_3bit_0/comp_p_3/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X74 uo_out[6] flashADC_3bit_0/comp_p_3/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X75 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_3/tail VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=20.433426 ps=144.985 w=10 l=1
X76 flashADC_3bit_0/comp_p_3/tail flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_3/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.5942 ps=82.28 w=9.995 l=0.35
X77 flashADC_3bit_0/comp_p_3/tail ua[0] flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.295525 ps=79.645 w=9.995 l=0.35
X78 flashADC_3bit_0/comp_p_3/tail ua[0] flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X79 flashADC_3bit_0/comp_p_3/tail ua[0] flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X80 flashADC_3bit_0/comp_p_3/tail ua[0] flashADC_3bit_0/comp_p_3/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X81 flashADC_3bit_0/comp_p_3/tail flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_3/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X82 flashADC_3bit_0/comp_p_3/tail flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_3/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X83 flashADC_3bit_0/comp_p_3/tail flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_3/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X84 flashADC_3bit_0/comp_p_4/latch_right flashADC_3bit_0/comp_p_4/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=5 l=1
X85 VDPWR flashADC_3bit_0/comp_p_4/out_left uo_out[7] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X86 flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/comp_p_4/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=4 l=1
X87 flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/comp_p_4/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=5 l=1
X88 flashADC_3bit_0/comp_p_4/latch_right flashADC_3bit_0/comp_p_4/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
X89 VDPWR flashADC_3bit_0/comp_p_4/out_left flashADC_3bit_0/comp_p_4/out_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X90 flashADC_3bit_0/comp_p_4/out_left flashADC_3bit_0/comp_p_4/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X91 uo_out[7] flashADC_3bit_0/comp_p_4/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X92 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_4/tail VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=20.433426 ps=144.985 w=10 l=1
X93 flashADC_3bit_0/comp_p_4/tail flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_4/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.5942 ps=82.28 w=9.995 l=0.35
X94 flashADC_3bit_0/comp_p_4/tail ua[0] flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.295525 ps=79.645 w=9.995 l=0.35
X95 flashADC_3bit_0/comp_p_4/tail ua[0] flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X96 flashADC_3bit_0/comp_p_4/tail ua[0] flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X97 flashADC_3bit_0/comp_p_4/tail ua[0] flashADC_3bit_0/comp_p_4/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X98 flashADC_3bit_0/comp_p_4/tail flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_4/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X99 flashADC_3bit_0/comp_p_4/tail flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_4/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X100 flashADC_3bit_0/comp_p_4/tail flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_4/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X101 flashADC_3bit_0/comp_p_5/latch_right flashADC_3bit_0/comp_p_5/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=5 l=1
X102 VDPWR flashADC_3bit_0/comp_p_5/out_left uio_out[0] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X103 flashADC_3bit_0/comp_p_5/latch_left flashADC_3bit_0/comp_p_5/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=4 l=1
X104 flashADC_3bit_0/comp_p_5/latch_left flashADC_3bit_0/comp_p_5/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=5 l=1
X105 flashADC_3bit_0/comp_p_5/latch_right flashADC_3bit_0/comp_p_5/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
X106 VDPWR flashADC_3bit_0/comp_p_5/out_left flashADC_3bit_0/comp_p_5/out_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X107 flashADC_3bit_0/comp_p_5/out_left flashADC_3bit_0/comp_p_5/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X108 uio_out[0] flashADC_3bit_0/comp_p_5/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X109 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_5/tail VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=20.433426 ps=144.985 w=10 l=1
X110 flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_5/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.5942 ps=82.28 w=9.995 l=0.35
X111 flashADC_3bit_0/comp_p_5/tail ua[0] flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.295525 ps=79.645 w=9.995 l=0.35
X112 flashADC_3bit_0/comp_p_5/tail ua[0] flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X113 flashADC_3bit_0/comp_p_5/tail ua[0] flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X114 flashADC_3bit_0/comp_p_5/tail ua[0] flashADC_3bit_0/comp_p_5/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X115 flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_5/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X116 flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_5/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X117 flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_5/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X118 flashADC_3bit_0/comp_p_6/latch_right flashADC_3bit_0/comp_p_6/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=5 l=1
X119 VDPWR flashADC_3bit_0/comp_p_6/out_left uio_out[1] VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X120 flashADC_3bit_0/comp_p_6/latch_left flashADC_3bit_0/comp_p_6/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=2.61 pd=19.16 as=0 ps=0 w=4 l=1
X121 flashADC_3bit_0/comp_p_6/latch_left flashADC_3bit_0/comp_p_6/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=5 l=1
X122 flashADC_3bit_0/comp_p_6/latch_right flashADC_3bit_0/comp_p_6/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
X123 VDPWR flashADC_3bit_0/comp_p_6/out_left flashADC_3bit_0/comp_p_6/out_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=1
X124 flashADC_3bit_0/comp_p_6/out_left flashADC_3bit_0/comp_p_6/latch_left VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X125 uio_out[1] flashADC_3bit_0/comp_p_6/latch_right VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=1
X126 VDPWR flashADC_3bit_0/comp_p_6/vbias_p flashADC_3bit_0/comp_p_6/tail VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=20.433426 ps=144.985 w=10 l=1
X127 flashADC_3bit_0/comp_p_6/tail flashADC_3bit_0/comp_p_6/vinn flashADC_3bit_0/comp_p_6/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.5942 ps=82.28 w=9.995 l=0.35
X128 flashADC_3bit_0/comp_p_6/tail ua[0] flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=11.295525 ps=79.645 w=9.995 l=0.35
X129 flashADC_3bit_0/comp_p_6/tail ua[0] flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X130 flashADC_3bit_0/comp_p_6/tail ua[0] flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X131 flashADC_3bit_0/comp_p_6/tail ua[0] flashADC_3bit_0/comp_p_6/latch_right VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X132 flashADC_3bit_0/comp_p_6/tail flashADC_3bit_0/comp_p_6/vinn flashADC_3bit_0/comp_p_6/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X133 flashADC_3bit_0/comp_p_6/tail flashADC_3bit_0/comp_p_6/vinn flashADC_3bit_0/comp_p_6/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X134 flashADC_3bit_0/comp_p_6/tail flashADC_3bit_0/comp_p_6/vinn flashADC_3bit_0/comp_p_6/latch_left VDPWR sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=9.995 l=0.35
X135 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X136 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X137 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out VDPWR sky130_fd_pr__pfet_01v8 ad=1.16 pd=9.16 as=1.16 ps=9.16 w=2 l=0.15
X138 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0.58 ps=5.16 w=1 l=0.15
X139 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VDPWR sky130_fd_pr__pfet_01v8 ad=1.16 pd=9.16 as=0 ps=0 w=2 l=0.15
X140 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X141 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X142 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X143 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out VDPWR sky130_fd_pr__pfet_01v8 ad=1.74 pd=13.74 as=1.16 ps=9.16 w=2 l=0.15
X144 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out VGND sky130_fd_pr__nfet_01v8 ad=0.87 pd=7.74 as=0.58 ps=5.16 w=1 l=0.15
X145 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B VDPWR sky130_fd_pr__pfet_01v8 ad=1.16 pd=9.16 as=0 ps=0 w=2 l=0.15
X146 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X147 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X148 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X149 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A VDPWR sky130_fd_pr__pfet_01v8 ad=1.16 pd=9.16 as=1.74 ps=13.74 w=2 l=0.15
X150 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0.87 ps=7.74 w=1 l=0.15
X151 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in VDPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
X152 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
R0 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 sky130_fd_pr__res_generic_m1 w=1 l=1
X153 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X154 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin uo_out[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X155 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X156 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=1.16 pd=9.16 as=0 ps=0 w=2 l=0.15
X157 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X158 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin uo_out[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X159 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X160 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_1/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
X161 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X162 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin uo_out[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X163 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X164 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_2/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
X165 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X166 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin uo_out[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X167 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X168 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R2 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_3/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X169 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X170 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin uo_out[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X171 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.15
X172 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=1.16 pd=9.16 as=0 ps=0 w=2 l=0.15
X173 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin uio_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X174 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin uio_out[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X175 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X176 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
X177 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin uio_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X178 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin uio_out[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X179 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X180 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
X181 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X182 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/in VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X183 uo_out[0] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X184 uo_out[0] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_7/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X185 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X186 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X187 uo_out[1] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X188 uo_out[1] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X189 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X190 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X191 uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X192 uo_out[2] flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_9/inv_1/vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X193 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X194 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X195 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out VDPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
X196 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_0/out VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X197 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A VDPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
X198 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
C0 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out 3.099387f
C1 flashADC_3bit_0/comp_p_6/vbias_p VDPWR 38.48766f
C2 flashADC_3bit_0/comp_p_1/latch_left flashADC_3bit_0/comp_p_1/tail 8.829929f
C3 ua[0] flashADC_3bit_0/comp_p_3/tail 2.919896f
C4 ua[0] flashADC_3bit_0/comp_p_4/tail 2.929377f
C5 uo_out[3] VDPWR 6.002129f
C6 ua[0] ua[1] 4.587688f
C7 uo_out[7] uio_out[0] 5.514357f
C8 uo_out[5] uo_out[4] 4.141313f
C9 flashADC_3bit_0/comp_p_1/latch_left flashADC_3bit_0/comp_p_1/latch_right 5.38251f
C10 flashADC_3bit_0/comp_p_4/out_left VDPWR 5.559441f
C11 uio_out[1] VDPWR 10.264361f
C12 flashADC_3bit_0/comp_p_0/tail flashADC_3bit_0/comp_p_0/latch_right 8.894202f
C13 flashADC_3bit_0/comp_p_2/tail flashADC_3bit_0/comp_p_2/latch_left 8.829929f
C14 flashADC_3bit_0/comp_p_1/vinn flashADC_3bit_0/comp_p_1/latch_right 3.543062f
C15 VDPWR uo_out[4] 4.888728f
C16 flashADC_3bit_0/comp_p_0/tail flashADC_3bit_0/comp_p_0/latch_left 8.829929f
C17 flashADC_3bit_0/comp_p_6/vinn VDPWR 3.827528f
C18 VDPWR flashADC_3bit_0/comp_p_5/out_left 7.450001f
C19 VDPWR flashADC_3bit_0/comp_p_6/latch_left 3.86486f
C20 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_6/out 5.14186f
C21 flashADC_3bit_0/comp_p_0/tail VDPWR 3.412349f
C22 flashADC_3bit_0/comp_p_2/out_left VDPWR 5.337812f
C23 flashADC_3bit_0/comp_p_3/latch_left VDPWR 3.721098f
C24 VDPWR flashADC_3bit_0/comp_p_1/tail 3.793449f
C25 flashADC_3bit_0/comp_p_4/vinn flashADC_3bit_0/comp_p_4/latch_right 3.536513f
C26 flashADC_3bit_0/comp_p_3/vinn flashADC_3bit_0/comp_p_3/latch_right 3.543126f
C27 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VDPWR 2.240643f
C28 VDPWR flashADC_3bit_0/comp_p_6/tail 3.765405f
C29 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_2/tail 8.894202f
C30 ua[0] flashADC_3bit_0/comp_p_6/vinn 2.274422f
C31 ua[0] flashADC_3bit_0/comp_p_0/tail 2.929379f
C32 VDPWR flashADC_3bit_0/comp_p_3/latch_right 3.668148f
C33 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_2/latch_left 5.38251f
C34 VDPWR flashADC_3bit_0/comp_p_1/latch_right 3.635097f
C35 uo_out[7] VDPWR 6.225174f
C36 flashADC_3bit_0/comp_p_0/out_left VDPWR 5.310384f
C37 flashADC_3bit_0/comp_p_6/vinn flashADC_3bit_0/comp_p_6/latch_right 3.538029f
C38 flashADC_3bit_0/comp_p_6/latch_left flashADC_3bit_0/comp_p_6/latch_right 5.38251f
C39 uio_out[0] VDPWR 6.487221f
C40 ua[0] flashADC_3bit_0/comp_p_1/tail 2.919898f
C41 flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/comp_p_4/latch_right 5.38251f
C42 flashADC_3bit_0/comp_p_3/latch_left flashADC_3bit_0/comp_p_3/tail 8.829929f
C43 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 5.877276f
C44 flashADC_3bit_0/comp_p_2/tail VDPWR 3.412596f
C45 flashADC_3bit_0/comp_p_0/vinn flashADC_3bit_0/comp_p_0/latch_right 3.537437f
C46 flashADC_3bit_0/comp_p_1/latch_left VDPWR 3.674756f
C47 ua[0] flashADC_3bit_0/comp_p_6/tail 2.917751f
C48 flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/comp_p_5/latch_right 8.894202f
C49 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out VDPWR 3.855608f
C50 flashADC_3bit_0/comp_p_1/out_left VDPWR 7.112554f
C51 flashADC_3bit_0/comp_p_6/latch_right flashADC_3bit_0/comp_p_6/tail 8.894202f
C52 flashADC_3bit_0/comp_p_5/latch_left flashADC_3bit_0/comp_p_5/latch_right 5.38251f
C53 flashADC_3bit_0/comp_p_1/vinn VDPWR 4.93284f
C54 flashADC_3bit_0/comp_p_3/tail flashADC_3bit_0/comp_p_3/latch_right 8.894202f
C55 uo_out[7] uo_out[6] 3.730491f
C56 VDPWR flashADC_3bit_0/comp_p_0/vinn 4.181973f
C57 flashADC_3bit_0/comp_p_4/latch_right flashADC_3bit_0/comp_p_4/tail 8.894202f
C58 VDPWR flashADC_3bit_0/comp_p_5/latch_right 3.785408f
C59 ua[0] flashADC_3bit_0/comp_p_2/tail 2.927971f
C60 flashADC_3bit_0/comp_p_5/vinn flashADC_3bit_0/comp_p_5/latch_right 3.543092f
C61 flashADC_3bit_0/comp_p_0/latch_left flashADC_3bit_0/comp_p_0/latch_right 5.38251f
C62 flashADC_3bit_0/comp_p_5/tail flashADC_3bit_0/comp_p_5/latch_left 8.829929f
C63 uo_out[5] VDPWR 5.495997f
C64 ua[0] flashADC_3bit_0/comp_p_1/vinn 2.227492f
C65 flashADC_3bit_0/comp_p_5/tail VDPWR 4.549301f
C66 ua[0] flashADC_3bit_0/comp_p_0/vinn 2.071417f
C67 flashADC_3bit_0/comp_p_3/vinn VDPWR 5.39465f
C68 flashADC_3bit_0/comp_p_4/vinn VDPWR 2.9131f
C69 VDPWR flashADC_3bit_0/comp_p_5/latch_left 3.828259f
C70 uo_out[5] uo_out[6] 3.339223f
C71 VDPWR flashADC_3bit_0/comp_p_6/out_left 7.102404f
C72 ua[0] flashADC_3bit_0/comp_p_5/tail 2.919896f
C73 VDPWR flashADC_3bit_0/comp_p_3/out_left 7.147648f
C74 VDPWR flashADC_3bit_0/comp_p_5/vinn 6.938992f
C75 uio_out[0] uio_out[1] 5.40212f
C76 flashADC_3bit_0/comp_p_6/latch_left flashADC_3bit_0/comp_p_6/tail 8.829929f
C77 ua[0] VDPWR 46.25895f
C78 VDPWR uo_out[6] 6.047353f
C79 VDPWR flashADC_3bit_0/comp_p_3/tail 3.799379f
C80 flashADC_3bit_0/comp_p_2/latch_right flashADC_3bit_0/comp_p_2/vinn 3.535519f
C81 VDPWR flashADC_3bit_0/comp_p_6/latch_right 3.794241f
C82 flashADC_3bit_0/comp_p_4/tail VDPWR 4.078566f
C83 VDPWR flashADC_3bit_0/tmux_7therm_to_3bin_0/tmux_2to1_3/B 2.389502f
C84 flashADC_3bit_0/comp_p_3/latch_left flashADC_3bit_0/comp_p_3/latch_right 5.38251f
C85 flashADC_3bit_0/comp_p_1/tail flashADC_3bit_0/comp_p_1/latch_right 8.894202f
C86 uo_out[1] uo_out[2] 2.072569f
C87 flashADC_3bit_0/comp_p_4/latch_left flashADC_3bit_0/comp_p_4/tail 8.829929f
C88 flashADC_3bit_0/comp_p_2/vinn VDPWR 2.400864f
C89 uo_out[2] VGND 2.349572f
C90 uio_out[1] VGND 7.953496f
C91 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_5/out VGND 2.050039f
C92 VDPWR VGND 0.491881p
C93 uio_out[0] VGND 6.02942f
C94 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_4/out VGND 2.162482f
C95 uo_out[7] VGND 12.596722f
C96 uo_out[6] VGND 5.369418f
C97 uo_out[5] VGND 9.80866f
C98 uo_out[4] VGND 9.897362f
C99 uo_out[3] VGND 5.921635f
C100 flashADC_3bit_0/tmux_7therm_to_3bin_0/buffer_8/in VGND 2.604635f
C101 flashADC_3bit_0/tmux_7therm_to_3bin_0/R1/R1 VGND 6.241027f
C102 ua[0] VGND 44.503277f
C103 flashADC_3bit_0/comp_p_6/vbias_p VGND 21.721624f
C104 flashADC_3bit_0/comp_p_6/latch_right VGND 5.891695f **FLOATING
C105 flashADC_3bit_0/comp_p_6/out_left VGND 3.852109f **FLOATING
C106 flashADC_3bit_0/comp_p_6/latch_left VGND 6.228204f **FLOATING
C107 flashADC_3bit_0/comp_p_5/latch_right VGND 5.563138f **FLOATING
C108 flashADC_3bit_0/comp_p_5/out_left VGND 3.765435f **FLOATING
C109 flashADC_3bit_0/comp_p_5/latch_left VGND 5.928939f **FLOATING
C110 flashADC_3bit_0/comp_p_4/latch_right VGND 7.574977f **FLOATING
C111 flashADC_3bit_0/comp_p_4/out_left VGND 6.007029f **FLOATING
C112 flashADC_3bit_0/comp_p_4/latch_left VGND 8.27735f **FLOATING
C113 flashADC_3bit_0/comp_p_3/latch_right VGND 5.619754f **FLOATING
C114 flashADC_3bit_0/comp_p_3/out_left VGND 4.205698f **FLOATING
C115 flashADC_3bit_0/comp_p_3/latch_left VGND 5.97815f **FLOATING
C116 flashADC_3bit_0/comp_p_2/latch_right VGND 7.590996f **FLOATING
C117 flashADC_3bit_0/comp_p_2/out_left VGND 6.327859f **FLOATING
C118 flashADC_3bit_0/comp_p_2/latch_left VGND 8.297646f **FLOATING
C119 flashADC_3bit_0/comp_p_0/latch_right VGND 7.581673f **FLOATING
C120 flashADC_3bit_0/comp_p_0/out_left VGND 6.310432f **FLOATING
C121 flashADC_3bit_0/comp_p_0/latch_left VGND 8.287999f **FLOATING
C122 flashADC_3bit_0/comp_p_1/latch_right VGND 5.574545f **FLOATING
C123 flashADC_3bit_0/comp_p_1/out_left VGND 4.11581f **FLOATING
C124 flashADC_3bit_0/comp_p_1/latch_left VGND 5.944707f **FLOATING
C125 flashADC_3bit_0/comp_p_1/vinn VGND 8.658644f
C126 flashADC_3bit_0/comp_p_0/vinn VGND 6.298379f
C127 flashADC_3bit_0/comp_p_2/vinn VGND 4.906179f
C128 flashADC_3bit_0/comp_p_3/vinn VGND 9.608513f
C129 flashADC_3bit_0/comp_p_4/vinn VGND 4.568718f
C130 flashADC_3bit_0/comp_p_5/vinn VGND 7.112859f
C131 flashADC_3bit_0/comp_p_6/vinn VGND 9.79437f
C132 ua[1] VGND 25.594332f
C133 flashADC_3bit_0/vbias_generation_0/bias_n VGND 3.404843f
C134 flashADC_3bit_0/vbias_generation_0/XR_bias_3/R2 VGND 2.006146f
